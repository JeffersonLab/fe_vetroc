LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY SRL16 IS
GENERIC
(
	INIT	: bit_vector := x"0000"
);
PORT
(
	Q		: OUT STD_LOGIC;
	A0		: IN STD_LOGIC;
	A1		: IN STD_LOGIC;
	A2		: IN STD_LOGIC;
	A3		: IN STD_LOGIC;
	CLK		: IN STD_LOGIC;
	D		: IN STD_LOGIC
);
END SRL16;

ARCHITECTURE srl16_arch OF SRL16 IS
	SIGNAL addr	: STD_LOGIC_VECTOR(3 DOWNTO 0);
	SIGNAL sr	: STD_LOGIC_VECTOR(15 DOWNTO 0) := x"0000";
BEGIN
	
	Q <= sr(CONV_INTEGER(addr));
	addr <= A3 & A2 & A1 & A0;

	PROCESS(CLK)
	BEGIN
		IF rising_edge(CLK) THEN
			sr <= sr(14 DOWNTO 0) & D;
		END IF;
	END PROCESS;
	
END srl16_arch;