-- megafunction wizard: %ALTGX_RECONFIG%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: alt2gxb_reconfig 

-- ============================================================
-- File Name: reconfig_side.vhd
-- Megafunction Name(s):
-- 			alt2gxb_reconfig
--
-- Simulation Library Files(s):
-- 			altera_mf;lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--alt2gxb_reconfig BASE_PORT_WIDTH=1 CBX_AUTO_BLACKBOX="ALL" CHANNEL_ADDRESS_WIDTH=8 DEVICE_FAMILY="Stratix IV" ENABLE_BUF_CAL="TRUE" ENABLE_CHL_ADDR_FOR_ANALOG_CTRL="TRUE" ENABLE_DFE="ON" ENABLE_EYE_MONITOR="ON" ENABLE_ILLEGAL_MODE_CHECK="TRUE" ENABLE_SELF_RECOVERY="TRUE" NUMBER_OF_CHANNELS=144 NUMBER_OF_RECONFIG_PORTS=36 READ_BASE_PORT_WIDTH=1 RECONFIG_FROMGXB_WIDTH=612 RECONFIG_MODE_SEL_WIDTH=4 RECONFIG_TOGXB_WIDTH=4 RX_EQDCGAIN_PORT_WIDTH=3 TX_PREEMP_PORT_WIDTH=5 busy ctrl_address ctrl_read ctrl_readdata ctrl_waitrequest ctrl_write ctrl_writedata data_valid error logical_channel_address read reconfig_clk reconfig_fromgxb reconfig_mode_sel reconfig_togxb rx_eqctrl rx_eqctrl_out rx_eqdcgain rx_eqdcgain_out tx_preemp_0t tx_preemp_0t_out tx_preemp_1t tx_preemp_1t_out tx_preemp_2t tx_preemp_2t_out tx_vodctrl tx_vodctrl_out write_all
--VERSION_BEGIN 13.0 cbx_alt2gxb_reconfig 2013:06:12:18:03:33:SJ cbx_alt_cal 2013:06:12:18:03:33:SJ cbx_alt_dprio 2013:06:12:18:03:33:SJ cbx_altsyncram 2013:06:12:18:03:33:SJ cbx_cycloneii 2013:06:12:18:03:33:SJ cbx_lpm_add_sub 2013:06:12:18:03:33:SJ cbx_lpm_compare 2013:06:12:18:03:33:SJ cbx_lpm_counter 2013:06:12:18:03:33:SJ cbx_lpm_decode 2013:06:12:18:03:33:SJ cbx_lpm_mux 2013:06:12:18:03:33:SJ cbx_lpm_shiftreg 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ cbx_stratix 2013:06:12:18:03:33:SJ cbx_stratixii 2013:06:12:18:03:33:SJ cbx_stratixiii 2013:06:12:18:03:33:SJ cbx_stratixv 2013:06:12:18:03:33:SJ cbx_util_mgl 2013:06:12:18:03:33:SJ  VERSION_END


--alt_dprio address_width=16 CBX_AUTO_BLACKBOX="ALL" device_family="Stratix IV" quad_address_width=9 address busy datain dataout dpclk dpriodisable dprioin dprioload dprioout quad_address rden reset wren wren_data
--VERSION_BEGIN 13.0 cbx_alt_dprio 2013:06:12:18:03:33:SJ cbx_cycloneii 2013:06:12:18:03:33:SJ cbx_lpm_add_sub 2013:06:12:18:03:33:SJ cbx_lpm_compare 2013:06:12:18:03:33:SJ cbx_lpm_counter 2013:06:12:18:03:33:SJ cbx_lpm_decode 2013:06:12:18:03:33:SJ cbx_lpm_shiftreg 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ cbx_stratix 2013:06:12:18:03:33:SJ cbx_stratixii 2013:06:12:18:03:33:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_compare 3 lpm_counter 1 lpm_decode 1 lut 1 reg 102 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  reconfig_side_alt_dprio_2vj IS 
	 PORT 
	 ( 
		 address	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 busy	:	OUT  STD_LOGIC;
		 datain	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
		 dataout	:	OUT  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 dpclk	:	IN  STD_LOGIC;
		 dpriodisable	:	OUT  STD_LOGIC;
		 dprioin	:	OUT  STD_LOGIC;
		 dprioload	:	OUT  STD_LOGIC;
		 dprioout	:	IN  STD_LOGIC;
		 quad_address	:	IN  STD_LOGIC_VECTOR (8 DOWNTO 0);
		 rden	:	IN  STD_LOGIC := '0';
		 reset	:	IN  STD_LOGIC := '0';
		 wren	:	IN  STD_LOGIC := '0';
		 wren_data	:	IN  STD_LOGIC := '0'
	 ); 
 END reconfig_side_alt_dprio_2vj;

 ARCHITECTURE RTL OF reconfig_side_alt_dprio_2vj IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "{-to addr_shift_reg[31]} DPRIO_INTERFACE_REG=ON;{-to wr_out_data_shift_reg[31]} DPRIO_INTERFACE_REG=ON;{-to rd_out_data_shift_reg[13]} DPRIO_INTERFACE_REG=ON;{-to in_data_shift_reg[0]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[0]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[1]} DPRIO_INTERFACE_REG=ON;{-to startup_cntr[2]} DPRIO_INTERFACE_REG=ON";

	 SIGNAL	 wire_addr_shift_reg_d	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wire_addr_shift_reg_asdata	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 addr_shift_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF addr_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_addr_shift_reg_w_q_range1337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 in_data_shift_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF in_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_rd_out_data_shift_reg_d	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL	 wire_rd_out_data_shift_reg_asdata	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL	 rd_out_data_shift_reg	:	STD_LOGIC_VECTOR(15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rd_out_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_rd_out_data_shift_reg_w_q_range1513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_startup_cntr_d	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL	 startup_cntr	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF startup_cntr : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_startup_cntr_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1578w1581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1582w1588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1582w1591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1574w1575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1574w1590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1574w1579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_lg_w_q_range1582w1583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range1574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range1578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_startup_cntr_w_q_range1582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 state_mc_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF state_mc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_state_mc_reg_w_q_range1172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range1191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range1207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_wr_out_data_shift_reg_d	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wire_wr_out_data_shift_reg_asdata	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL	 wr_out_data_shift_reg	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_out_data_shift_reg : SIGNAL IS "PRESERVE_REGISTER=ON;POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_wr_out_data_shift_reg_w_q_range1448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_w_lg_agb1335w1512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_w_lg_agb1335w1447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_w_lg_agb1335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_pre_amble_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_pre_amble_cmpr_agb	:	STD_LOGIC;
	 SIGNAL  wire_pre_amble_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_rd_data_output_cmpr_ageb	:	STD_LOGIC;
	 SIGNAL  wire_rd_data_output_cmpr_alb	:	STD_LOGIC;
	 SIGNAL  wire_rd_data_output_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_cmpr_aeb	:	STD_LOGIC;
	 SIGNAL  wire_state_mc_cmpr_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_counter_cnt_en	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_write_state1157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_counter_q	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_state_mc_decode_eq	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL	wire_dprioin_mux_dataout	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s0_to_01174w1175w1176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s1_to_01193w1194w1195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_s2_to_01209w1210w1211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wren1163w1186w1199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wren1163w1186w1187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_wr_addr_state1334w1338w1339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rd_data_output_state1514w1515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wr_data_state1449w1450w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s0_to_01174w1175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s1_to_01193w1194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_s2_to_01209w1210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren1163w1186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren1163w1164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wren1163w1181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_w_lg_rden1570w1571w1572w1573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_wr_addr_state1334w1338w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state1200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state1182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state1189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state1166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_idle_state1203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rd_data_output_state1514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wr_data_state1449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_01174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_11173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_01193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_11192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_01209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_11208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_startup_done1568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_startup_idle1569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren1163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren_data1185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_rden1570w1571w1572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rden1161w1162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_rden1570w1571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rden1161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rden1570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rdinc1198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_rdinc1180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s0_to_11177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s1_to_11196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_s2_to_11212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wr_addr_state1334w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren1188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren1165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_wren1202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  busy_state :	STD_LOGIC;
	 SIGNAL  idle_state :	STD_LOGIC;
	 SIGNAL  rd_addr_done :	STD_LOGIC;
	 SIGNAL  rd_addr_state :	STD_LOGIC;
	 SIGNAL  rd_data_done :	STD_LOGIC;
	 SIGNAL  rd_data_input_state :	STD_LOGIC;
	 SIGNAL  rd_data_output_state :	STD_LOGIC;
	 SIGNAL  rd_data_state :	STD_LOGIC;
	 SIGNAL  rdinc	:	STD_LOGIC;
	 SIGNAL  read_state :	STD_LOGIC;
	 SIGNAL  s0_to_0 :	STD_LOGIC;
	 SIGNAL  s0_to_1 :	STD_LOGIC;
	 SIGNAL  s1_to_0 :	STD_LOGIC;
	 SIGNAL  s1_to_1 :	STD_LOGIC;
	 SIGNAL  s2_to_0 :	STD_LOGIC;
	 SIGNAL  s2_to_1 :	STD_LOGIC;
	 SIGNAL  startup_done :	STD_LOGIC;
	 SIGNAL  startup_idle :	STD_LOGIC;
	 SIGNAL  wr_addr_done :	STD_LOGIC;
	 SIGNAL  wr_addr_state :	STD_LOGIC;
	 SIGNAL  wr_data_done :	STD_LOGIC;
	 SIGNAL  wr_data_state :	STD_LOGIC;
	 SIGNAL  write_state :	STD_LOGIC;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_decode
	 GENERIC 
	 (
		LPM_DECODES	:	NATURAL;
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_decode"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		enable	:	IN STD_LOGIC := '1';
		eq	:	OUT STD_LOGIC_VECTOR(LPM_DECODES-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_dprio_w_lg_w_lg_w_lg_s0_to_01174w1175w1176w(0) <= wire_dprio_w_lg_w_lg_s0_to_01174w1175w(0) AND wire_state_mc_reg_w_q_range1172w(0);
	wire_dprio_w_lg_w_lg_w_lg_s1_to_01193w1194w1195w(0) <= wire_dprio_w_lg_w_lg_s1_to_01193w1194w(0) AND wire_state_mc_reg_w_q_range1191w(0);
	wire_dprio_w_lg_w_lg_w_lg_s2_to_01209w1210w1211w(0) <= wire_dprio_w_lg_w_lg_s2_to_01209w1210w(0) AND wire_state_mc_reg_w_q_range1207w(0);
	wire_dprio_w_lg_w_lg_w_lg_wren1163w1186w1199w(0) <= wire_dprio_w_lg_w_lg_wren1163w1186w(0) AND wire_dprio_w_lg_rdinc1198w(0);
	wire_dprio_w_lg_w_lg_w_lg_wren1163w1186w1187w(0) <= wire_dprio_w_lg_w_lg_wren1163w1186w(0) AND rden;
	wire_dprio_w_lg_w_lg_w_lg_wr_addr_state1334w1338w1339w(0) <= wire_dprio_w_lg_w_lg_wr_addr_state1334w1338w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_rd_data_output_state1514w1515w(0) <= wire_dprio_w_lg_rd_data_output_state1514w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_wr_data_state1449w1450w(0) <= wire_dprio_w_lg_wr_data_state1449w(0) AND wire_pre_amble_cmpr_agb;
	wire_dprio_w_lg_w_lg_s0_to_01174w1175w(0) <= wire_dprio_w_lg_s0_to_01174w(0) AND wire_dprio_w_lg_s0_to_11173w(0);
	wire_dprio_w_lg_w_lg_s1_to_01193w1194w(0) <= wire_dprio_w_lg_s1_to_01193w(0) AND wire_dprio_w_lg_s1_to_11192w(0);
	wire_dprio_w_lg_w_lg_s2_to_01209w1210w(0) <= wire_dprio_w_lg_s2_to_01209w(0) AND wire_dprio_w_lg_s2_to_11208w(0);
	wire_dprio_w_lg_w_lg_wren1163w1186w(0) <= wire_dprio_w_lg_wren1163w(0) AND wire_dprio_w_lg_wren_data1185w(0);
	wire_dprio_w_lg_w_lg_wren1163w1164w(0) <= wire_dprio_w_lg_wren1163w(0) AND wire_dprio_w_lg_w_lg_rden1161w1162w(0);
	wire_dprio_w_lg_w_lg_wren1163w1181w(0) <= wire_dprio_w_lg_wren1163w(0) AND wire_dprio_w_lg_rdinc1180w(0);
	wire_dprio_w_lg_w_lg_w_lg_w_lg_rden1570w1571w1572w1573w(0) <= wire_dprio_w_lg_w_lg_w_lg_rden1570w1571w1572w(0) AND wire_dprio_w_lg_startup_done1568w(0);
	wire_dprio_w_lg_w_lg_wr_addr_state1334w1338w(0) <= wire_dprio_w_lg_wr_addr_state1334w(0) AND wire_addr_shift_reg_w_q_range1337w(0);
	wire_dprio_w_lg_idle_state1200w(0) <= idle_state AND wire_dprio_w_lg_w_lg_w_lg_wren1163w1186w1199w(0);
	wire_dprio_w_lg_idle_state1182w(0) <= idle_state AND wire_dprio_w_lg_w_lg_wren1163w1181w(0);
	wire_dprio_w_lg_idle_state1189w(0) <= idle_state AND wire_dprio_w_lg_wren1188w(0);
	wire_dprio_w_lg_idle_state1166w(0) <= idle_state AND wire_dprio_w_lg_wren1165w(0);
	wire_dprio_w_lg_idle_state1203w(0) <= idle_state AND wire_dprio_w_lg_wren1202w(0);
	wire_dprio_w_lg_rd_data_output_state1514w(0) <= rd_data_output_state AND wire_rd_out_data_shift_reg_w_q_range1513w(0);
	wire_dprio_w_lg_wr_data_state1449w(0) <= wr_data_state AND wire_wr_out_data_shift_reg_w_q_range1448w(0);
	wire_dprio_w_lg_s0_to_01174w(0) <= NOT s0_to_0;
	wire_dprio_w_lg_s0_to_11173w(0) <= NOT s0_to_1;
	wire_dprio_w_lg_s1_to_01193w(0) <= NOT s1_to_0;
	wire_dprio_w_lg_s1_to_11192w(0) <= NOT s1_to_1;
	wire_dprio_w_lg_s2_to_01209w(0) <= NOT s2_to_0;
	wire_dprio_w_lg_s2_to_11208w(0) <= NOT s2_to_1;
	wire_dprio_w_lg_startup_done1568w(0) <= NOT startup_done;
	wire_dprio_w_lg_startup_idle1569w(0) <= NOT startup_idle;
	wire_dprio_w_lg_wren1163w(0) <= NOT wren;
	wire_dprio_w_lg_wren_data1185w(0) <= NOT wren_data;
	wire_dprio_w_lg_w_lg_w_lg_rden1570w1571w1572w(0) <= wire_dprio_w_lg_w_lg_rden1570w1571w(0) OR wire_dprio_w_lg_startup_idle1569w(0);
	wire_dprio_w_lg_w_lg_rden1161w1162w(0) <= wire_dprio_w_lg_rden1161w(0) OR wren_data;
	wire_dprio_w_lg_w_lg_rden1570w1571w(0) <= wire_dprio_w_lg_rden1570w(0) OR rdinc;
	wire_dprio_w_lg_rden1161w(0) <= rden OR rdinc;
	wire_dprio_w_lg_rden1570w(0) <= rden OR wren;
	wire_dprio_w_lg_rdinc1198w(0) <= rdinc OR rden;
	wire_dprio_w_lg_rdinc1180w(0) <= rdinc OR wren_data;
	wire_dprio_w_lg_s0_to_11177w(0) <= s0_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s0_to_01174w1175w1176w(0);
	wire_dprio_w_lg_s1_to_11196w(0) <= s1_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s1_to_01193w1194w1195w(0);
	wire_dprio_w_lg_s2_to_11212w(0) <= s2_to_1 OR wire_dprio_w_lg_w_lg_w_lg_s2_to_01209w1210w1211w(0);
	wire_dprio_w_lg_wr_addr_state1334w(0) <= wr_addr_state OR rd_addr_state;
	wire_dprio_w_lg_wren1188w(0) <= wren OR wire_dprio_w_lg_w_lg_w_lg_wren1163w1186w1187w(0);
	wire_dprio_w_lg_wren1165w(0) <= wren OR wire_dprio_w_lg_w_lg_wren1163w1164w(0);
	wire_dprio_w_lg_wren1202w(0) <= wren OR wren_data;
	busy <= busy_state;
	busy_state <= (write_state OR read_state);
	dataout <= in_data_shift_reg;
	dpriodisable <= (NOT wire_startup_cntr_w_lg_w_q_range1582w1591w(0));
	dprioin <= wire_dprioin_mux_dataout;
	dprioload <= (NOT (wire_startup_cntr_w_lg_w_q_range1574w1579w(0) AND (NOT startup_cntr(2))));
	idle_state <= wire_state_mc_decode_eq(0);
	rd_addr_done <= (rd_addr_state AND wire_state_mc_cmpr_aeb);
	rd_addr_state <= (wire_state_mc_decode_eq(5) AND startup_done);
	rd_data_done <= (rd_data_state AND wire_state_mc_cmpr_aeb);
	rd_data_input_state <= (wire_rd_data_output_cmpr_ageb AND rd_data_state);
	rd_data_output_state <= (wire_rd_data_output_cmpr_alb AND rd_data_state);
	rd_data_state <= (wire_state_mc_decode_eq(7) AND startup_done);
	rdinc <= '0';
	read_state <= (rd_addr_state OR rd_data_state);
	s0_to_0 <= ((wr_data_state AND wr_data_done) OR (rd_data_state AND rd_data_done));
	s0_to_1 <= ((wire_dprio_w_lg_idle_state1166w(0) OR (wr_addr_state AND wr_addr_done)) OR (rd_addr_state AND rd_addr_done));
	s1_to_0 <= (((wr_data_state AND wr_data_done) OR (rd_data_state AND rd_data_done)) OR wire_dprio_w_lg_idle_state1189w(0));
	s1_to_1 <= ((wire_dprio_w_lg_idle_state1182w(0) OR (wr_addr_state AND wr_addr_done)) OR (rd_addr_state AND rd_addr_done));
	s2_to_0 <= ((((wr_addr_state AND wr_addr_done) OR (wr_data_state AND wr_data_done)) OR (rd_data_state AND rd_data_done)) OR wire_dprio_w_lg_idle_state1203w(0));
	s2_to_1 <= (wire_dprio_w_lg_idle_state1200w(0) OR (rd_addr_state AND rd_addr_done));
	startup_done <= (wire_startup_cntr_w_lg_w_q_range1582w1588w(0) AND startup_cntr(1));
	startup_idle <= (wire_startup_cntr_w_lg_w_q_range1574w1575w(0) AND (NOT (startup_cntr(2) XOR startup_cntr(1))));
	wr_addr_done <= (wr_addr_state AND wire_state_mc_cmpr_aeb);
	wr_addr_state <= (wire_state_mc_decode_eq(1) AND startup_done);
	wr_data_done <= (wr_data_state AND wire_state_mc_cmpr_aeb);
	wr_data_state <= (wire_state_mc_decode_eq(3) AND startup_done);
	write_state <= (wr_addr_state OR wr_data_state);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(0) <= wire_addr_shift_reg_asdata(0);
				ELSE addr_shift_reg(0) <= wire_addr_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(1) <= wire_addr_shift_reg_asdata(1);
				ELSE addr_shift_reg(1) <= wire_addr_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(2) <= wire_addr_shift_reg_asdata(2);
				ELSE addr_shift_reg(2) <= wire_addr_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(3) <= wire_addr_shift_reg_asdata(3);
				ELSE addr_shift_reg(3) <= wire_addr_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(4) <= wire_addr_shift_reg_asdata(4);
				ELSE addr_shift_reg(4) <= wire_addr_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(5) <= wire_addr_shift_reg_asdata(5);
				ELSE addr_shift_reg(5) <= wire_addr_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(6) <= wire_addr_shift_reg_asdata(6);
				ELSE addr_shift_reg(6) <= wire_addr_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(7) <= wire_addr_shift_reg_asdata(7);
				ELSE addr_shift_reg(7) <= wire_addr_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(8) <= wire_addr_shift_reg_asdata(8);
				ELSE addr_shift_reg(8) <= wire_addr_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(9) <= wire_addr_shift_reg_asdata(9);
				ELSE addr_shift_reg(9) <= wire_addr_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(10) <= wire_addr_shift_reg_asdata(10);
				ELSE addr_shift_reg(10) <= wire_addr_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(11) <= wire_addr_shift_reg_asdata(11);
				ELSE addr_shift_reg(11) <= wire_addr_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(12) <= wire_addr_shift_reg_asdata(12);
				ELSE addr_shift_reg(12) <= wire_addr_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(13) <= wire_addr_shift_reg_asdata(13);
				ELSE addr_shift_reg(13) <= wire_addr_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(14) <= wire_addr_shift_reg_asdata(14);
				ELSE addr_shift_reg(14) <= wire_addr_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(15) <= wire_addr_shift_reg_asdata(15);
				ELSE addr_shift_reg(15) <= wire_addr_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(16) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(16) <= wire_addr_shift_reg_asdata(16);
				ELSE addr_shift_reg(16) <= wire_addr_shift_reg_d(16);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(17) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(17) <= wire_addr_shift_reg_asdata(17);
				ELSE addr_shift_reg(17) <= wire_addr_shift_reg_d(17);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(18) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(18) <= wire_addr_shift_reg_asdata(18);
				ELSE addr_shift_reg(18) <= wire_addr_shift_reg_d(18);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(19) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(19) <= wire_addr_shift_reg_asdata(19);
				ELSE addr_shift_reg(19) <= wire_addr_shift_reg_d(19);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(20) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(20) <= wire_addr_shift_reg_asdata(20);
				ELSE addr_shift_reg(20) <= wire_addr_shift_reg_d(20);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(21) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(21) <= wire_addr_shift_reg_asdata(21);
				ELSE addr_shift_reg(21) <= wire_addr_shift_reg_d(21);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(22) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(22) <= wire_addr_shift_reg_asdata(22);
				ELSE addr_shift_reg(22) <= wire_addr_shift_reg_d(22);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(23) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(23) <= wire_addr_shift_reg_asdata(23);
				ELSE addr_shift_reg(23) <= wire_addr_shift_reg_d(23);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(24) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(24) <= wire_addr_shift_reg_asdata(24);
				ELSE addr_shift_reg(24) <= wire_addr_shift_reg_d(24);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(25) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(25) <= wire_addr_shift_reg_asdata(25);
				ELSE addr_shift_reg(25) <= wire_addr_shift_reg_d(25);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(26) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(26) <= wire_addr_shift_reg_asdata(26);
				ELSE addr_shift_reg(26) <= wire_addr_shift_reg_d(26);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(27) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(27) <= wire_addr_shift_reg_asdata(27);
				ELSE addr_shift_reg(27) <= wire_addr_shift_reg_d(27);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(28) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(28) <= wire_addr_shift_reg_asdata(28);
				ELSE addr_shift_reg(28) <= wire_addr_shift_reg_d(28);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(29) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(29) <= wire_addr_shift_reg_asdata(29);
				ELSE addr_shift_reg(29) <= wire_addr_shift_reg_d(29);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(30) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(30) <= wire_addr_shift_reg_asdata(30);
				ELSE addr_shift_reg(30) <= wire_addr_shift_reg_d(30);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN addr_shift_reg(31) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN addr_shift_reg(31) <= wire_addr_shift_reg_asdata(31);
				ELSE addr_shift_reg(31) <= wire_addr_shift_reg_d(31);
				END IF;
		END IF;
	END PROCESS;
	wire_addr_shift_reg_asdata <= ( "00" & "00" & "0" & quad_address(8 DOWNTO 0) & "10" & address);
	wire_addr_shift_reg_d <= ( addr_shift_reg(30 DOWNTO 0) & "0");
	wire_addr_shift_reg_w_q_range1337w(0) <= addr_shift_reg(31);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN in_data_shift_reg <= (OTHERS => '0');
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
			IF (rd_data_input_state = '1') THEN in_data_shift_reg <= ( in_data_shift_reg(14 DOWNTO 0) & dprioout);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(0) <= wire_rd_out_data_shift_reg_asdata(0);
				ELSE rd_out_data_shift_reg(0) <= wire_rd_out_data_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(1) <= wire_rd_out_data_shift_reg_asdata(1);
				ELSE rd_out_data_shift_reg(1) <= wire_rd_out_data_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(2) <= wire_rd_out_data_shift_reg_asdata(2);
				ELSE rd_out_data_shift_reg(2) <= wire_rd_out_data_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(3) <= wire_rd_out_data_shift_reg_asdata(3);
				ELSE rd_out_data_shift_reg(3) <= wire_rd_out_data_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(4) <= wire_rd_out_data_shift_reg_asdata(4);
				ELSE rd_out_data_shift_reg(4) <= wire_rd_out_data_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(5) <= wire_rd_out_data_shift_reg_asdata(5);
				ELSE rd_out_data_shift_reg(5) <= wire_rd_out_data_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(6) <= wire_rd_out_data_shift_reg_asdata(6);
				ELSE rd_out_data_shift_reg(6) <= wire_rd_out_data_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(7) <= wire_rd_out_data_shift_reg_asdata(7);
				ELSE rd_out_data_shift_reg(7) <= wire_rd_out_data_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(8) <= wire_rd_out_data_shift_reg_asdata(8);
				ELSE rd_out_data_shift_reg(8) <= wire_rd_out_data_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(9) <= wire_rd_out_data_shift_reg_asdata(9);
				ELSE rd_out_data_shift_reg(9) <= wire_rd_out_data_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(10) <= wire_rd_out_data_shift_reg_asdata(10);
				ELSE rd_out_data_shift_reg(10) <= wire_rd_out_data_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(11) <= wire_rd_out_data_shift_reg_asdata(11);
				ELSE rd_out_data_shift_reg(11) <= wire_rd_out_data_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(12) <= wire_rd_out_data_shift_reg_asdata(12);
				ELSE rd_out_data_shift_reg(12) <= wire_rd_out_data_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(13) <= wire_rd_out_data_shift_reg_asdata(13);
				ELSE rd_out_data_shift_reg(13) <= wire_rd_out_data_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(14) <= wire_rd_out_data_shift_reg_asdata(14);
				ELSE rd_out_data_shift_reg(14) <= wire_rd_out_data_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN rd_out_data_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN rd_out_data_shift_reg(15) <= wire_rd_out_data_shift_reg_asdata(15);
				ELSE rd_out_data_shift_reg(15) <= wire_rd_out_data_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	wire_rd_out_data_shift_reg_asdata <= ( "00" & "1" & "1" & "0" & quad_address & "10");
	wire_rd_out_data_shift_reg_d <= ( rd_out_data_shift_reg(14 DOWNTO 0) & "0");
	wire_rd_out_data_shift_reg_w_q_range1513w(0) <= rd_out_data_shift_reg(15);
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(0) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(0) <= '0';
				ELSE startup_cntr(0) <= wire_startup_cntr_d(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(1) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(1) <= '0';
				ELSE startup_cntr(1) <= wire_startup_cntr_d(1);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk)
	BEGIN
		IF (dpclk = '1' AND dpclk'event) THEN 
			IF (wire_startup_cntr_ena(2) = '1') THEN 
				IF (reset = '1') THEN startup_cntr(2) <= '0';
				ELSE startup_cntr(2) <= wire_startup_cntr_d(2);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_startup_cntr_d <= ( wire_startup_cntr_w_lg_w_q_range1582w1583w & wire_startup_cntr_w_lg_w_q_range1574w1579w & wire_startup_cntr_w_lg_w_q_range1574w1575w);
	loop0 : FOR i IN 0 TO 2 GENERATE
		wire_startup_cntr_ena(i) <= wire_dprio_w_lg_w_lg_w_lg_w_lg_rden1570w1571w1572w1573w(0);
	END GENERATE loop0;
	wire_startup_cntr_w_lg_w_q_range1578w1581w(0) <= wire_startup_cntr_w_q_range1578w(0) AND wire_startup_cntr_w_q_range1574w(0);
	wire_startup_cntr_w_lg_w_q_range1582w1588w(0) <= wire_startup_cntr_w_q_range1582w(0) AND wire_startup_cntr_w_lg_w_q_range1574w1575w(0);
	wire_startup_cntr_w_lg_w_q_range1582w1591w(0) <= wire_startup_cntr_w_q_range1582w(0) AND wire_startup_cntr_w_lg_w_q_range1574w1590w(0);
	wire_startup_cntr_w_lg_w_q_range1574w1575w(0) <= NOT wire_startup_cntr_w_q_range1574w(0);
	wire_startup_cntr_w_lg_w_q_range1574w1590w(0) <= wire_startup_cntr_w_q_range1574w(0) OR wire_startup_cntr_w_q_range1578w(0);
	wire_startup_cntr_w_lg_w_q_range1574w1579w(0) <= wire_startup_cntr_w_q_range1574w(0) XOR wire_startup_cntr_w_q_range1578w(0);
	wire_startup_cntr_w_lg_w_q_range1582w1583w(0) <= wire_startup_cntr_w_q_range1582w(0) XOR wire_startup_cntr_w_lg_w_q_range1578w1581w(0);
	wire_startup_cntr_w_q_range1574w(0) <= startup_cntr(0);
	wire_startup_cntr_w_q_range1578w(0) <= startup_cntr(1);
	wire_startup_cntr_w_q_range1582w(0) <= startup_cntr(2);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN state_mc_reg <= (OTHERS => '0');
		ELSIF (dpclk = '1' AND dpclk'event) THEN state_mc_reg <= ( wire_dprio_w_lg_s2_to_11212w & wire_dprio_w_lg_s1_to_11196w & wire_dprio_w_lg_s0_to_11177w);
		END IF;
	END PROCESS;
	wire_state_mc_reg_w_q_range1172w(0) <= state_mc_reg(0);
	wire_state_mc_reg_w_q_range1191w(0) <= state_mc_reg(1);
	wire_state_mc_reg_w_q_range1207w(0) <= state_mc_reg(2);
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(0) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(0) <= wire_wr_out_data_shift_reg_asdata(0);
				ELSE wr_out_data_shift_reg(0) <= wire_wr_out_data_shift_reg_d(0);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(1) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(1) <= wire_wr_out_data_shift_reg_asdata(1);
				ELSE wr_out_data_shift_reg(1) <= wire_wr_out_data_shift_reg_d(1);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(2) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(2) <= wire_wr_out_data_shift_reg_asdata(2);
				ELSE wr_out_data_shift_reg(2) <= wire_wr_out_data_shift_reg_d(2);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(3) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(3) <= wire_wr_out_data_shift_reg_asdata(3);
				ELSE wr_out_data_shift_reg(3) <= wire_wr_out_data_shift_reg_d(3);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(4) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(4) <= wire_wr_out_data_shift_reg_asdata(4);
				ELSE wr_out_data_shift_reg(4) <= wire_wr_out_data_shift_reg_d(4);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(5) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(5) <= wire_wr_out_data_shift_reg_asdata(5);
				ELSE wr_out_data_shift_reg(5) <= wire_wr_out_data_shift_reg_d(5);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(6) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(6) <= wire_wr_out_data_shift_reg_asdata(6);
				ELSE wr_out_data_shift_reg(6) <= wire_wr_out_data_shift_reg_d(6);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(7) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(7) <= wire_wr_out_data_shift_reg_asdata(7);
				ELSE wr_out_data_shift_reg(7) <= wire_wr_out_data_shift_reg_d(7);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(8) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(8) <= wire_wr_out_data_shift_reg_asdata(8);
				ELSE wr_out_data_shift_reg(8) <= wire_wr_out_data_shift_reg_d(8);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(9) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(9) <= wire_wr_out_data_shift_reg_asdata(9);
				ELSE wr_out_data_shift_reg(9) <= wire_wr_out_data_shift_reg_d(9);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(10) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(10) <= wire_wr_out_data_shift_reg_asdata(10);
				ELSE wr_out_data_shift_reg(10) <= wire_wr_out_data_shift_reg_d(10);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(11) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(11) <= wire_wr_out_data_shift_reg_asdata(11);
				ELSE wr_out_data_shift_reg(11) <= wire_wr_out_data_shift_reg_d(11);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(12) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(12) <= wire_wr_out_data_shift_reg_asdata(12);
				ELSE wr_out_data_shift_reg(12) <= wire_wr_out_data_shift_reg_d(12);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(13) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(13) <= wire_wr_out_data_shift_reg_asdata(13);
				ELSE wr_out_data_shift_reg(13) <= wire_wr_out_data_shift_reg_d(13);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(14) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(14) <= wire_wr_out_data_shift_reg_asdata(14);
				ELSE wr_out_data_shift_reg(14) <= wire_wr_out_data_shift_reg_d(14);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(15) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(15) <= wire_wr_out_data_shift_reg_asdata(15);
				ELSE wr_out_data_shift_reg(15) <= wire_wr_out_data_shift_reg_d(15);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(16) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(16) <= wire_wr_out_data_shift_reg_asdata(16);
				ELSE wr_out_data_shift_reg(16) <= wire_wr_out_data_shift_reg_d(16);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(17) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(17) <= wire_wr_out_data_shift_reg_asdata(17);
				ELSE wr_out_data_shift_reg(17) <= wire_wr_out_data_shift_reg_d(17);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(18) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(18) <= wire_wr_out_data_shift_reg_asdata(18);
				ELSE wr_out_data_shift_reg(18) <= wire_wr_out_data_shift_reg_d(18);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(19) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(19) <= wire_wr_out_data_shift_reg_asdata(19);
				ELSE wr_out_data_shift_reg(19) <= wire_wr_out_data_shift_reg_d(19);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(20) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(20) <= wire_wr_out_data_shift_reg_asdata(20);
				ELSE wr_out_data_shift_reg(20) <= wire_wr_out_data_shift_reg_d(20);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(21) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(21) <= wire_wr_out_data_shift_reg_asdata(21);
				ELSE wr_out_data_shift_reg(21) <= wire_wr_out_data_shift_reg_d(21);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(22) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(22) <= wire_wr_out_data_shift_reg_asdata(22);
				ELSE wr_out_data_shift_reg(22) <= wire_wr_out_data_shift_reg_d(22);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(23) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(23) <= wire_wr_out_data_shift_reg_asdata(23);
				ELSE wr_out_data_shift_reg(23) <= wire_wr_out_data_shift_reg_d(23);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(24) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(24) <= wire_wr_out_data_shift_reg_asdata(24);
				ELSE wr_out_data_shift_reg(24) <= wire_wr_out_data_shift_reg_d(24);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(25) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(25) <= wire_wr_out_data_shift_reg_asdata(25);
				ELSE wr_out_data_shift_reg(25) <= wire_wr_out_data_shift_reg_d(25);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(26) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(26) <= wire_wr_out_data_shift_reg_asdata(26);
				ELSE wr_out_data_shift_reg(26) <= wire_wr_out_data_shift_reg_d(26);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(27) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(27) <= wire_wr_out_data_shift_reg_asdata(27);
				ELSE wr_out_data_shift_reg(27) <= wire_wr_out_data_shift_reg_d(27);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(28) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(28) <= wire_wr_out_data_shift_reg_asdata(28);
				ELSE wr_out_data_shift_reg(28) <= wire_wr_out_data_shift_reg_d(28);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(29) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(29) <= wire_wr_out_data_shift_reg_asdata(29);
				ELSE wr_out_data_shift_reg(29) <= wire_wr_out_data_shift_reg_d(29);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(30) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(30) <= wire_wr_out_data_shift_reg_asdata(30);
				ELSE wr_out_data_shift_reg(30) <= wire_wr_out_data_shift_reg_d(30);
				END IF;
		END IF;
	END PROCESS;
	PROCESS (dpclk, reset)
	BEGIN
		IF (reset = '1') THEN wr_out_data_shift_reg(31) <= '0';
		ELSIF (dpclk = '1' AND dpclk'event) THEN 
				IF (wire_pre_amble_cmpr_aeb = '1') THEN wr_out_data_shift_reg(31) <= wire_wr_out_data_shift_reg_asdata(31);
				ELSE wr_out_data_shift_reg(31) <= wire_wr_out_data_shift_reg_d(31);
				END IF;
		END IF;
	END PROCESS;
	wire_wr_out_data_shift_reg_asdata <= ( "00" & "01" & "0" & quad_address(8 DOWNTO 0) & "10" & datain);
	wire_wr_out_data_shift_reg_d <= ( wr_out_data_shift_reg(30 DOWNTO 0) & "0");
	wire_wr_out_data_shift_reg_w_q_range1448w(0) <= wr_out_data_shift_reg(31);
	wire_pre_amble_cmpr_w_lg_w_lg_agb1335w1512w(0) <= wire_pre_amble_cmpr_w_lg_agb1335w(0) AND rd_data_output_state;
	wire_pre_amble_cmpr_w_lg_w_lg_agb1335w1447w(0) <= wire_pre_amble_cmpr_w_lg_agb1335w(0) AND wr_data_state;
	wire_pre_amble_cmpr_w_lg_agb1335w(0) <= NOT wire_pre_amble_cmpr_agb;
	wire_pre_amble_cmpr_datab <= "011111";
	pre_amble_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_pre_amble_cmpr_aeb,
		agb => wire_pre_amble_cmpr_agb,
		dataa => wire_state_mc_counter_q,
		datab => wire_pre_amble_cmpr_datab
	  );
	wire_rd_data_output_cmpr_datab <= "110000";
	rd_data_output_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		ageb => wire_rd_data_output_cmpr_ageb,
		alb => wire_rd_data_output_cmpr_alb,
		dataa => wire_state_mc_counter_q,
		datab => wire_rd_data_output_cmpr_datab
	  );
	wire_state_mc_cmpr_datab <= (OTHERS => '1');
	state_mc_cmpr :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		aeb => wire_state_mc_cmpr_aeb,
		dataa => wire_state_mc_counter_q,
		datab => wire_state_mc_cmpr_datab
	  );
	wire_state_mc_counter_cnt_en <= wire_dprio_w_lg_write_state1157w(0);
	wire_dprio_w_lg_write_state1157w(0) <= write_state OR read_state;
	state_mc_counter :  lpm_counter
	  GENERIC MAP (
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 6
	  )
	  PORT MAP ( 
		clock => dpclk,
		cnt_en => wire_state_mc_counter_cnt_en,
		q => wire_state_mc_counter_q,
		sclr => reset
	  );
	state_mc_decode :  lpm_decode
	  GENERIC MAP (
		LPM_DECODES => 8,
		LPM_WIDTH => 3
	  )
	  PORT MAP ( 
		data => state_mc_reg,
		eq => wire_state_mc_decode_eq
	  );
	wire_dprioin_mux_dataout <= (((wire_dprio_w_lg_w_lg_w_lg_wr_addr_state1334w1338w1339w(0) OR (wire_pre_amble_cmpr_w_lg_agb1335w(0) AND wire_dprio_w_lg_wr_addr_state1334w(0))) OR (wire_dprio_w_lg_w_lg_wr_data_state1449w1450w(0) OR wire_pre_amble_cmpr_w_lg_w_lg_agb1335w1447w(0))) OR (wire_dprio_w_lg_w_lg_rd_data_output_state1514w1515w(0) OR wire_pre_amble_cmpr_w_lg_w_lg_agb1335w1512w(0))) OR NOT(((write_state OR rd_addr_state) OR rd_data_output_state));

 END RTL; --reconfig_side_alt_dprio_2vj


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" LPM_SIZE=4 LPM_WIDTH=16 LPM_WIDTHS=2 data result sel
--VERSION_BEGIN 13.0 cbx_lpm_mux 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ  VERSION_END

--synthesis_resources = lut 16 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  reconfig_side_mux_t7a IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END reconfig_side_mux_t7a;

 ARCHITECTURE RTL OF reconfig_side_mux_t7a IS

	 SIGNAL	wire_l1_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w10_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w10_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w11_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w11_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w12_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w12_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w13_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w13_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w14_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w14_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w15_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w15_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w5_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w5_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w6_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w6_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w7_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w7_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w8_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w8_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w9_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w9_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w10_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w11_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w12_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w13_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w14_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w15_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w1_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w2_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w3_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w4_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w5_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w6_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w7_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w8_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w9_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL  data_wire :	STD_LOGIC_VECTOR (95 DOWNTO 0);
	 SIGNAL  result_wire_ext :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  sel_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
 BEGIN

	data_wire <= ( wire_l1_w15_n1_mux_dataout & wire_l1_w15_n0_mux_dataout & wire_l1_w14_n1_mux_dataout & wire_l1_w14_n0_mux_dataout & wire_l1_w13_n1_mux_dataout & wire_l1_w13_n0_mux_dataout & wire_l1_w12_n1_mux_dataout & wire_l1_w12_n0_mux_dataout & wire_l1_w11_n1_mux_dataout & wire_l1_w11_n0_mux_dataout & wire_l1_w10_n1_mux_dataout & wire_l1_w10_n0_mux_dataout & wire_l1_w9_n1_mux_dataout & wire_l1_w9_n0_mux_dataout & wire_l1_w8_n1_mux_dataout & wire_l1_w8_n0_mux_dataout & wire_l1_w7_n1_mux_dataout & wire_l1_w7_n0_mux_dataout & wire_l1_w6_n1_mux_dataout & wire_l1_w6_n0_mux_dataout & wire_l1_w5_n1_mux_dataout & wire_l1_w5_n0_mux_dataout & wire_l1_w4_n1_mux_dataout & wire_l1_w4_n0_mux_dataout & wire_l1_w3_n1_mux_dataout & wire_l1_w3_n0_mux_dataout & wire_l1_w2_n1_mux_dataout & wire_l1_w2_n0_mux_dataout & wire_l1_w1_n1_mux_dataout & wire_l1_w1_n0_mux_dataout & wire_l1_w0_n1_mux_dataout & wire_l1_w0_n0_mux_dataout & data);
	result <= result_wire_ext;
	result_wire_ext <= ( wire_l2_w15_n0_mux_dataout & wire_l2_w14_n0_mux_dataout & wire_l2_w13_n0_mux_dataout & wire_l2_w12_n0_mux_dataout & wire_l2_w11_n0_mux_dataout & wire_l2_w10_n0_mux_dataout & wire_l2_w9_n0_mux_dataout & wire_l2_w8_n0_mux_dataout & wire_l2_w7_n0_mux_dataout & wire_l2_w6_n0_mux_dataout & wire_l2_w5_n0_mux_dataout & wire_l2_w4_n0_mux_dataout & wire_l2_w3_n0_mux_dataout & wire_l2_w2_n0_mux_dataout & wire_l2_w1_n0_mux_dataout & wire_l2_w0_n0_mux_dataout);
	sel_wire <= ( sel(1) & "00" & sel(0));
	wire_l1_w0_n0_mux_dataout <= data_wire(16) WHEN sel_wire(0) = '1'  ELSE data_wire(0);
	wire_l1_w0_n1_mux_dataout <= data_wire(48) WHEN sel_wire(0) = '1'  ELSE data_wire(32);
	wire_l1_w10_n0_mux_dataout <= data_wire(26) WHEN sel_wire(0) = '1'  ELSE data_wire(10);
	wire_l1_w10_n1_mux_dataout <= data_wire(58) WHEN sel_wire(0) = '1'  ELSE data_wire(42);
	wire_l1_w11_n0_mux_dataout <= data_wire(27) WHEN sel_wire(0) = '1'  ELSE data_wire(11);
	wire_l1_w11_n1_mux_dataout <= data_wire(59) WHEN sel_wire(0) = '1'  ELSE data_wire(43);
	wire_l1_w12_n0_mux_dataout <= data_wire(28) WHEN sel_wire(0) = '1'  ELSE data_wire(12);
	wire_l1_w12_n1_mux_dataout <= data_wire(60) WHEN sel_wire(0) = '1'  ELSE data_wire(44);
	wire_l1_w13_n0_mux_dataout <= data_wire(29) WHEN sel_wire(0) = '1'  ELSE data_wire(13);
	wire_l1_w13_n1_mux_dataout <= data_wire(61) WHEN sel_wire(0) = '1'  ELSE data_wire(45);
	wire_l1_w14_n0_mux_dataout <= data_wire(30) WHEN sel_wire(0) = '1'  ELSE data_wire(14);
	wire_l1_w14_n1_mux_dataout <= data_wire(62) WHEN sel_wire(0) = '1'  ELSE data_wire(46);
	wire_l1_w15_n0_mux_dataout <= data_wire(31) WHEN sel_wire(0) = '1'  ELSE data_wire(15);
	wire_l1_w15_n1_mux_dataout <= data_wire(63) WHEN sel_wire(0) = '1'  ELSE data_wire(47);
	wire_l1_w1_n0_mux_dataout <= data_wire(17) WHEN sel_wire(0) = '1'  ELSE data_wire(1);
	wire_l1_w1_n1_mux_dataout <= data_wire(49) WHEN sel_wire(0) = '1'  ELSE data_wire(33);
	wire_l1_w2_n0_mux_dataout <= data_wire(18) WHEN sel_wire(0) = '1'  ELSE data_wire(2);
	wire_l1_w2_n1_mux_dataout <= data_wire(50) WHEN sel_wire(0) = '1'  ELSE data_wire(34);
	wire_l1_w3_n0_mux_dataout <= data_wire(19) WHEN sel_wire(0) = '1'  ELSE data_wire(3);
	wire_l1_w3_n1_mux_dataout <= data_wire(51) WHEN sel_wire(0) = '1'  ELSE data_wire(35);
	wire_l1_w4_n0_mux_dataout <= data_wire(20) WHEN sel_wire(0) = '1'  ELSE data_wire(4);
	wire_l1_w4_n1_mux_dataout <= data_wire(52) WHEN sel_wire(0) = '1'  ELSE data_wire(36);
	wire_l1_w5_n0_mux_dataout <= data_wire(21) WHEN sel_wire(0) = '1'  ELSE data_wire(5);
	wire_l1_w5_n1_mux_dataout <= data_wire(53) WHEN sel_wire(0) = '1'  ELSE data_wire(37);
	wire_l1_w6_n0_mux_dataout <= data_wire(22) WHEN sel_wire(0) = '1'  ELSE data_wire(6);
	wire_l1_w6_n1_mux_dataout <= data_wire(54) WHEN sel_wire(0) = '1'  ELSE data_wire(38);
	wire_l1_w7_n0_mux_dataout <= data_wire(23) WHEN sel_wire(0) = '1'  ELSE data_wire(7);
	wire_l1_w7_n1_mux_dataout <= data_wire(55) WHEN sel_wire(0) = '1'  ELSE data_wire(39);
	wire_l1_w8_n0_mux_dataout <= data_wire(24) WHEN sel_wire(0) = '1'  ELSE data_wire(8);
	wire_l1_w8_n1_mux_dataout <= data_wire(56) WHEN sel_wire(0) = '1'  ELSE data_wire(40);
	wire_l1_w9_n0_mux_dataout <= data_wire(25) WHEN sel_wire(0) = '1'  ELSE data_wire(9);
	wire_l1_w9_n1_mux_dataout <= data_wire(57) WHEN sel_wire(0) = '1'  ELSE data_wire(41);
	wire_l2_w0_n0_mux_dataout <= data_wire(65) WHEN sel_wire(3) = '1'  ELSE data_wire(64);
	wire_l2_w10_n0_mux_dataout <= data_wire(85) WHEN sel_wire(3) = '1'  ELSE data_wire(84);
	wire_l2_w11_n0_mux_dataout <= data_wire(87) WHEN sel_wire(3) = '1'  ELSE data_wire(86);
	wire_l2_w12_n0_mux_dataout <= data_wire(89) WHEN sel_wire(3) = '1'  ELSE data_wire(88);
	wire_l2_w13_n0_mux_dataout <= data_wire(91) WHEN sel_wire(3) = '1'  ELSE data_wire(90);
	wire_l2_w14_n0_mux_dataout <= data_wire(93) WHEN sel_wire(3) = '1'  ELSE data_wire(92);
	wire_l2_w15_n0_mux_dataout <= data_wire(95) WHEN sel_wire(3) = '1'  ELSE data_wire(94);
	wire_l2_w1_n0_mux_dataout <= data_wire(67) WHEN sel_wire(3) = '1'  ELSE data_wire(66);
	wire_l2_w2_n0_mux_dataout <= data_wire(69) WHEN sel_wire(3) = '1'  ELSE data_wire(68);
	wire_l2_w3_n0_mux_dataout <= data_wire(71) WHEN sel_wire(3) = '1'  ELSE data_wire(70);
	wire_l2_w4_n0_mux_dataout <= data_wire(73) WHEN sel_wire(3) = '1'  ELSE data_wire(72);
	wire_l2_w5_n0_mux_dataout <= data_wire(75) WHEN sel_wire(3) = '1'  ELSE data_wire(74);
	wire_l2_w6_n0_mux_dataout <= data_wire(77) WHEN sel_wire(3) = '1'  ELSE data_wire(76);
	wire_l2_w7_n0_mux_dataout <= data_wire(79) WHEN sel_wire(3) = '1'  ELSE data_wire(78);
	wire_l2_w8_n0_mux_dataout <= data_wire(81) WHEN sel_wire(3) = '1'  ELSE data_wire(80);
	wire_l2_w9_n0_mux_dataout <= data_wire(83) WHEN sel_wire(3) = '1'  ELSE data_wire(82);

 END RTL; --reconfig_side_mux_t7a


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" LPM_SIZE=4 LPM_WIDTH=2 LPM_WIDTHS=2 data result sel
--VERSION_BEGIN 13.0 cbx_lpm_mux 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ  VERSION_END

--synthesis_resources = lut 2 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  reconfig_side_mux_86a IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (1 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END reconfig_side_mux_86a;

 ARCHITECTURE RTL OF reconfig_side_mux_86a IS

	 SIGNAL	wire_l1_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w1_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL  data_wire :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  result_wire_ext :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  sel_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
 BEGIN

	data_wire <= ( wire_l1_w1_n1_mux_dataout & wire_l1_w1_n0_mux_dataout & wire_l1_w0_n1_mux_dataout & wire_l1_w0_n0_mux_dataout & data);
	result <= result_wire_ext;
	result_wire_ext <= ( wire_l2_w1_n0_mux_dataout & wire_l2_w0_n0_mux_dataout);
	sel_wire <= ( sel(1) & "00" & sel(0));
	wire_l1_w0_n0_mux_dataout <= data_wire(2) WHEN sel_wire(0) = '1'  ELSE data_wire(0);
	wire_l1_w0_n1_mux_dataout <= data_wire(6) WHEN sel_wire(0) = '1'  ELSE data_wire(4);
	wire_l1_w1_n0_mux_dataout <= data_wire(3) WHEN sel_wire(0) = '1'  ELSE data_wire(1);
	wire_l1_w1_n1_mux_dataout <= data_wire(7) WHEN sel_wire(0) = '1'  ELSE data_wire(5);
	wire_l2_w0_n0_mux_dataout <= data_wire(9) WHEN sel_wire(3) = '1'  ELSE data_wire(8);
	wire_l2_w1_n0_mux_dataout <= data_wire(11) WHEN sel_wire(3) = '1'  ELSE data_wire(10);

 END RTL; --reconfig_side_mux_86a


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" LPM_SIZE=4 LPM_WIDTH=12 LPM_WIDTHS=2 data result sel
--VERSION_BEGIN 13.0 cbx_lpm_mux 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ  VERSION_END

--synthesis_resources = lut 12 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  reconfig_side_mux_p7a IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (47 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (11 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END reconfig_side_mux_p7a;

 ARCHITECTURE RTL OF reconfig_side_mux_p7a IS

	 SIGNAL	wire_l1_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w10_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w10_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w11_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w11_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w1_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w2_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w3_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w4_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w5_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w5_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w6_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w6_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w7_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w7_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w8_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w8_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w9_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w9_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w10_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w11_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w1_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w2_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w3_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w4_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w5_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w6_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w7_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w8_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w9_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL  data_wire :	STD_LOGIC_VECTOR (71 DOWNTO 0);
	 SIGNAL  result_wire_ext :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  sel_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
 BEGIN

	data_wire <= ( wire_l1_w11_n1_mux_dataout & wire_l1_w11_n0_mux_dataout & wire_l1_w10_n1_mux_dataout & wire_l1_w10_n0_mux_dataout & wire_l1_w9_n1_mux_dataout & wire_l1_w9_n0_mux_dataout & wire_l1_w8_n1_mux_dataout & wire_l1_w8_n0_mux_dataout & wire_l1_w7_n1_mux_dataout & wire_l1_w7_n0_mux_dataout & wire_l1_w6_n1_mux_dataout & wire_l1_w6_n0_mux_dataout & wire_l1_w5_n1_mux_dataout & wire_l1_w5_n0_mux_dataout & wire_l1_w4_n1_mux_dataout & wire_l1_w4_n0_mux_dataout & wire_l1_w3_n1_mux_dataout & wire_l1_w3_n0_mux_dataout & wire_l1_w2_n1_mux_dataout & wire_l1_w2_n0_mux_dataout & wire_l1_w1_n1_mux_dataout & wire_l1_w1_n0_mux_dataout & wire_l1_w0_n1_mux_dataout & wire_l1_w0_n0_mux_dataout & data);
	result <= result_wire_ext;
	result_wire_ext <= ( wire_l2_w11_n0_mux_dataout & wire_l2_w10_n0_mux_dataout & wire_l2_w9_n0_mux_dataout & wire_l2_w8_n0_mux_dataout & wire_l2_w7_n0_mux_dataout & wire_l2_w6_n0_mux_dataout & wire_l2_w5_n0_mux_dataout & wire_l2_w4_n0_mux_dataout & wire_l2_w3_n0_mux_dataout & wire_l2_w2_n0_mux_dataout & wire_l2_w1_n0_mux_dataout & wire_l2_w0_n0_mux_dataout);
	sel_wire <= ( sel(1) & "00" & sel(0));
	wire_l1_w0_n0_mux_dataout <= data_wire(12) WHEN sel_wire(0) = '1'  ELSE data_wire(0);
	wire_l1_w0_n1_mux_dataout <= data_wire(36) WHEN sel_wire(0) = '1'  ELSE data_wire(24);
	wire_l1_w10_n0_mux_dataout <= data_wire(22) WHEN sel_wire(0) = '1'  ELSE data_wire(10);
	wire_l1_w10_n1_mux_dataout <= data_wire(46) WHEN sel_wire(0) = '1'  ELSE data_wire(34);
	wire_l1_w11_n0_mux_dataout <= data_wire(23) WHEN sel_wire(0) = '1'  ELSE data_wire(11);
	wire_l1_w11_n1_mux_dataout <= data_wire(47) WHEN sel_wire(0) = '1'  ELSE data_wire(35);
	wire_l1_w1_n0_mux_dataout <= data_wire(13) WHEN sel_wire(0) = '1'  ELSE data_wire(1);
	wire_l1_w1_n1_mux_dataout <= data_wire(37) WHEN sel_wire(0) = '1'  ELSE data_wire(25);
	wire_l1_w2_n0_mux_dataout <= data_wire(14) WHEN sel_wire(0) = '1'  ELSE data_wire(2);
	wire_l1_w2_n1_mux_dataout <= data_wire(38) WHEN sel_wire(0) = '1'  ELSE data_wire(26);
	wire_l1_w3_n0_mux_dataout <= data_wire(15) WHEN sel_wire(0) = '1'  ELSE data_wire(3);
	wire_l1_w3_n1_mux_dataout <= data_wire(39) WHEN sel_wire(0) = '1'  ELSE data_wire(27);
	wire_l1_w4_n0_mux_dataout <= data_wire(16) WHEN sel_wire(0) = '1'  ELSE data_wire(4);
	wire_l1_w4_n1_mux_dataout <= data_wire(40) WHEN sel_wire(0) = '1'  ELSE data_wire(28);
	wire_l1_w5_n0_mux_dataout <= data_wire(17) WHEN sel_wire(0) = '1'  ELSE data_wire(5);
	wire_l1_w5_n1_mux_dataout <= data_wire(41) WHEN sel_wire(0) = '1'  ELSE data_wire(29);
	wire_l1_w6_n0_mux_dataout <= data_wire(18) WHEN sel_wire(0) = '1'  ELSE data_wire(6);
	wire_l1_w6_n1_mux_dataout <= data_wire(42) WHEN sel_wire(0) = '1'  ELSE data_wire(30);
	wire_l1_w7_n0_mux_dataout <= data_wire(19) WHEN sel_wire(0) = '1'  ELSE data_wire(7);
	wire_l1_w7_n1_mux_dataout <= data_wire(43) WHEN sel_wire(0) = '1'  ELSE data_wire(31);
	wire_l1_w8_n0_mux_dataout <= data_wire(20) WHEN sel_wire(0) = '1'  ELSE data_wire(8);
	wire_l1_w8_n1_mux_dataout <= data_wire(44) WHEN sel_wire(0) = '1'  ELSE data_wire(32);
	wire_l1_w9_n0_mux_dataout <= data_wire(21) WHEN sel_wire(0) = '1'  ELSE data_wire(9);
	wire_l1_w9_n1_mux_dataout <= data_wire(45) WHEN sel_wire(0) = '1'  ELSE data_wire(33);
	wire_l2_w0_n0_mux_dataout <= data_wire(49) WHEN sel_wire(3) = '1'  ELSE data_wire(48);
	wire_l2_w10_n0_mux_dataout <= data_wire(69) WHEN sel_wire(3) = '1'  ELSE data_wire(68);
	wire_l2_w11_n0_mux_dataout <= data_wire(71) WHEN sel_wire(3) = '1'  ELSE data_wire(70);
	wire_l2_w1_n0_mux_dataout <= data_wire(51) WHEN sel_wire(3) = '1'  ELSE data_wire(50);
	wire_l2_w2_n0_mux_dataout <= data_wire(53) WHEN sel_wire(3) = '1'  ELSE data_wire(52);
	wire_l2_w3_n0_mux_dataout <= data_wire(55) WHEN sel_wire(3) = '1'  ELSE data_wire(54);
	wire_l2_w4_n0_mux_dataout <= data_wire(57) WHEN sel_wire(3) = '1'  ELSE data_wire(56);
	wire_l2_w5_n0_mux_dataout <= data_wire(59) WHEN sel_wire(3) = '1'  ELSE data_wire(58);
	wire_l2_w6_n0_mux_dataout <= data_wire(61) WHEN sel_wire(3) = '1'  ELSE data_wire(60);
	wire_l2_w7_n0_mux_dataout <= data_wire(63) WHEN sel_wire(3) = '1'  ELSE data_wire(62);
	wire_l2_w8_n0_mux_dataout <= data_wire(65) WHEN sel_wire(3) = '1'  ELSE data_wire(64);
	wire_l2_w9_n0_mux_dataout <= data_wire(67) WHEN sel_wire(3) = '1'  ELSE data_wire(66);

 END RTL; --reconfig_side_mux_p7a


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" LPM_SIZE=144 LPM_WIDTH=1 LPM_WIDTHS=8 data result sel
--VERSION_BEGIN 13.0 cbx_lpm_mux 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ  VERSION_END

--synthesis_resources = lut 85 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  reconfig_side_mux_i9a IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (143 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END reconfig_side_mux_i9a;

 ARCHITECTURE RTL OF reconfig_side_mux_i9a IS

	 SIGNAL	wire_l1_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n100_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n101_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n102_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n103_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n104_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n105_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n106_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n107_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n108_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n109_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n10_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n110_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n111_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n112_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n113_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n114_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n115_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n116_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n117_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n118_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n119_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n11_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n120_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n121_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n122_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n123_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n124_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n125_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n126_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n127_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n12_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n13_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n14_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n15_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n16_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n17_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n18_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n19_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n20_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n21_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n22_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n23_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n24_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n25_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n26_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n27_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n28_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n29_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n30_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n31_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n32_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n33_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n34_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n35_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n36_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n37_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n38_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n39_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n40_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n41_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n42_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n43_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n44_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n45_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n46_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n47_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n48_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n49_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n4_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n50_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n51_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n52_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n53_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n54_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n55_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n56_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n57_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n58_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n59_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n5_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n60_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n61_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n62_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n63_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n64_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n65_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n66_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n67_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n68_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n69_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n6_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n70_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n71_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n72_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n73_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n74_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n75_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n76_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n77_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n78_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n79_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n7_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n80_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n81_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n82_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n83_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n84_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n85_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n86_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n87_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n88_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n89_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n8_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n90_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n91_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n92_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n93_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n94_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n95_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n96_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n97_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n98_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n99_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n9_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n10_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n11_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n12_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n13_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n14_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n15_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n16_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n17_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n18_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n19_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n20_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n21_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n22_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n23_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n24_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n25_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n26_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n27_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n28_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n29_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n30_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n31_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n32_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n33_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n34_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n35_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n36_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n37_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n38_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n39_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n40_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n41_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n42_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n43_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n44_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n45_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n46_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n47_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n48_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n49_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n4_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n50_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n51_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n52_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n53_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n54_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n55_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n56_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n57_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n58_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n59_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n5_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n60_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n61_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n62_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n63_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n6_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n7_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n8_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n9_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n10_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n11_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n12_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n13_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n14_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n15_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n16_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n17_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n18_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n19_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n20_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n21_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n22_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n23_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n24_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n25_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n26_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n27_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n28_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n29_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n30_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n31_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n4_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n5_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n6_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n7_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n8_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n9_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n10_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n11_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n12_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n13_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n14_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n15_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n4_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n5_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n6_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n7_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n8_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n9_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l5_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l5_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l5_w0_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l5_w0_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l5_w0_n4_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l5_w0_n5_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l5_w0_n6_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l5_w0_n7_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l6_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l6_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l6_w0_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l6_w0_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l7_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l7_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l8_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL  data_wire :	STD_LOGIC_VECTOR (509 DOWNTO 0);
	 SIGNAL  result_wire_ext :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  sel_wire :	STD_LOGIC_VECTOR (63 DOWNTO 0);
 BEGIN

	data_wire <= ( wire_l7_w0_n1_mux_dataout & wire_l7_w0_n0_mux_dataout & wire_l6_w0_n3_mux_dataout & wire_l6_w0_n2_mux_dataout & wire_l6_w0_n1_mux_dataout & wire_l6_w0_n0_mux_dataout & wire_l5_w0_n7_mux_dataout & wire_l5_w0_n6_mux_dataout & wire_l5_w0_n5_mux_dataout & wire_l5_w0_n4_mux_dataout & wire_l5_w0_n3_mux_dataout & wire_l5_w0_n2_mux_dataout & wire_l5_w0_n1_mux_dataout & wire_l5_w0_n0_mux_dataout & wire_l4_w0_n15_mux_dataout & wire_l4_w0_n14_mux_dataout & wire_l4_w0_n13_mux_dataout & wire_l4_w0_n12_mux_dataout & wire_l4_w0_n11_mux_dataout & wire_l4_w0_n10_mux_dataout & wire_l4_w0_n9_mux_dataout & wire_l4_w0_n8_mux_dataout & wire_l4_w0_n7_mux_dataout & wire_l4_w0_n6_mux_dataout & wire_l4_w0_n5_mux_dataout & wire_l4_w0_n4_mux_dataout & wire_l4_w0_n3_mux_dataout & wire_l4_w0_n2_mux_dataout & wire_l4_w0_n1_mux_dataout & wire_l4_w0_n0_mux_dataout & wire_l3_w0_n31_mux_dataout & wire_l3_w0_n30_mux_dataout & wire_l3_w0_n29_mux_dataout & wire_l3_w0_n28_mux_dataout & wire_l3_w0_n27_mux_dataout & wire_l3_w0_n26_mux_dataout & wire_l3_w0_n25_mux_dataout & wire_l3_w0_n24_mux_dataout & wire_l3_w0_n23_mux_dataout & wire_l3_w0_n22_mux_dataout & wire_l3_w0_n21_mux_dataout & wire_l3_w0_n20_mux_dataout & wire_l3_w0_n19_mux_dataout & wire_l3_w0_n18_mux_dataout & wire_l3_w0_n17_mux_dataout & wire_l3_w0_n16_mux_dataout & wire_l3_w0_n15_mux_dataout & wire_l3_w0_n14_mux_dataout & wire_l3_w0_n13_mux_dataout & wire_l3_w0_n12_mux_dataout & wire_l3_w0_n11_mux_dataout & wire_l3_w0_n10_mux_dataout & wire_l3_w0_n9_mux_dataout & wire_l3_w0_n8_mux_dataout & wire_l3_w0_n7_mux_dataout & wire_l3_w0_n6_mux_dataout & wire_l3_w0_n5_mux_dataout & wire_l3_w0_n4_mux_dataout & wire_l3_w0_n3_mux_dataout & wire_l3_w0_n2_mux_dataout & wire_l3_w0_n1_mux_dataout & wire_l3_w0_n0_mux_dataout & wire_l2_w0_n63_mux_dataout & wire_l2_w0_n62_mux_dataout & wire_l2_w0_n61_mux_dataout & wire_l2_w0_n60_mux_dataout & wire_l2_w0_n59_mux_dataout & wire_l2_w0_n58_mux_dataout & wire_l2_w0_n57_mux_dataout & wire_l2_w0_n56_mux_dataout & wire_l2_w0_n55_mux_dataout & wire_l2_w0_n54_mux_dataout
 & wire_l2_w0_n53_mux_dataout & wire_l2_w0_n52_mux_dataout & wire_l2_w0_n51_mux_dataout & wire_l2_w0_n50_mux_dataout & wire_l2_w0_n49_mux_dataout & wire_l2_w0_n48_mux_dataout & wire_l2_w0_n47_mux_dataout & wire_l2_w0_n46_mux_dataout & wire_l2_w0_n45_mux_dataout & wire_l2_w0_n44_mux_dataout & wire_l2_w0_n43_mux_dataout & wire_l2_w0_n42_mux_dataout & wire_l2_w0_n41_mux_dataout & wire_l2_w0_n40_mux_dataout & wire_l2_w0_n39_mux_dataout & wire_l2_w0_n38_mux_dataout & wire_l2_w0_n37_mux_dataout & wire_l2_w0_n36_mux_dataout & wire_l2_w0_n35_mux_dataout & wire_l2_w0_n34_mux_dataout & wire_l2_w0_n33_mux_dataout & wire_l2_w0_n32_mux_dataout & wire_l2_w0_n31_mux_dataout & wire_l2_w0_n30_mux_dataout & wire_l2_w0_n29_mux_dataout & wire_l2_w0_n28_mux_dataout & wire_l2_w0_n27_mux_dataout & wire_l2_w0_n26_mux_dataout & wire_l2_w0_n25_mux_dataout & wire_l2_w0_n24_mux_dataout & wire_l2_w0_n23_mux_dataout & wire_l2_w0_n22_mux_dataout & wire_l2_w0_n21_mux_dataout & wire_l2_w0_n20_mux_dataout & wire_l2_w0_n19_mux_dataout & wire_l2_w0_n18_mux_dataout & wire_l2_w0_n17_mux_dataout & wire_l2_w0_n16_mux_dataout & wire_l2_w0_n15_mux_dataout & wire_l2_w0_n14_mux_dataout & wire_l2_w0_n13_mux_dataout & wire_l2_w0_n12_mux_dataout & wire_l2_w0_n11_mux_dataout & wire_l2_w0_n10_mux_dataout & wire_l2_w0_n9_mux_dataout & wire_l2_w0_n8_mux_dataout & wire_l2_w0_n7_mux_dataout & wire_l2_w0_n6_mux_dataout & wire_l2_w0_n5_mux_dataout & wire_l2_w0_n4_mux_dataout & wire_l2_w0_n3_mux_dataout & wire_l2_w0_n2_mux_dataout & wire_l2_w0_n1_mux_dataout & wire_l2_w0_n0_mux_dataout & wire_l1_w0_n127_mux_dataout & wire_l1_w0_n126_mux_dataout & wire_l1_w0_n125_mux_dataout & wire_l1_w0_n124_mux_dataout & wire_l1_w0_n123_mux_dataout & wire_l1_w0_n122_mux_dataout & wire_l1_w0_n121_mux_dataout & wire_l1_w0_n120_mux_dataout & wire_l1_w0_n119_mux_dataout & wire_l1_w0_n118_mux_dataout & wire_l1_w0_n117_mux_dataout & wire_l1_w0_n116_mux_dataout & wire_l1_w0_n115_mux_dataout & wire_l1_w0_n114_mux_dataout & wire_l1_w0_n113_mux_dataout & wire_l1_w0_n112_mux_dataout & wire_l1_w0_n111_mux_dataout
 & wire_l1_w0_n110_mux_dataout & wire_l1_w0_n109_mux_dataout & wire_l1_w0_n108_mux_dataout & wire_l1_w0_n107_mux_dataout & wire_l1_w0_n106_mux_dataout & wire_l1_w0_n105_mux_dataout & wire_l1_w0_n104_mux_dataout & wire_l1_w0_n103_mux_dataout & wire_l1_w0_n102_mux_dataout & wire_l1_w0_n101_mux_dataout & wire_l1_w0_n100_mux_dataout & wire_l1_w0_n99_mux_dataout & wire_l1_w0_n98_mux_dataout & wire_l1_w0_n97_mux_dataout & wire_l1_w0_n96_mux_dataout & wire_l1_w0_n95_mux_dataout & wire_l1_w0_n94_mux_dataout & wire_l1_w0_n93_mux_dataout & wire_l1_w0_n92_mux_dataout & wire_l1_w0_n91_mux_dataout & wire_l1_w0_n90_mux_dataout & wire_l1_w0_n89_mux_dataout & wire_l1_w0_n88_mux_dataout & wire_l1_w0_n87_mux_dataout & wire_l1_w0_n86_mux_dataout & wire_l1_w0_n85_mux_dataout & wire_l1_w0_n84_mux_dataout & wire_l1_w0_n83_mux_dataout & wire_l1_w0_n82_mux_dataout & wire_l1_w0_n81_mux_dataout & wire_l1_w0_n80_mux_dataout & wire_l1_w0_n79_mux_dataout & wire_l1_w0_n78_mux_dataout & wire_l1_w0_n77_mux_dataout & wire_l1_w0_n76_mux_dataout & wire_l1_w0_n75_mux_dataout & wire_l1_w0_n74_mux_dataout & wire_l1_w0_n73_mux_dataout & wire_l1_w0_n72_mux_dataout & wire_l1_w0_n71_mux_dataout & wire_l1_w0_n70_mux_dataout & wire_l1_w0_n69_mux_dataout & wire_l1_w0_n68_mux_dataout & wire_l1_w0_n67_mux_dataout & wire_l1_w0_n66_mux_dataout & wire_l1_w0_n65_mux_dataout & wire_l1_w0_n64_mux_dataout & wire_l1_w0_n63_mux_dataout & wire_l1_w0_n62_mux_dataout & wire_l1_w0_n61_mux_dataout & wire_l1_w0_n60_mux_dataout & wire_l1_w0_n59_mux_dataout & wire_l1_w0_n58_mux_dataout & wire_l1_w0_n57_mux_dataout & wire_l1_w0_n56_mux_dataout & wire_l1_w0_n55_mux_dataout & wire_l1_w0_n54_mux_dataout & wire_l1_w0_n53_mux_dataout & wire_l1_w0_n52_mux_dataout & wire_l1_w0_n51_mux_dataout & wire_l1_w0_n50_mux_dataout & wire_l1_w0_n49_mux_dataout & wire_l1_w0_n48_mux_dataout & wire_l1_w0_n47_mux_dataout & wire_l1_w0_n46_mux_dataout & wire_l1_w0_n45_mux_dataout & wire_l1_w0_n44_mux_dataout & wire_l1_w0_n43_mux_dataout & wire_l1_w0_n42_mux_dataout & wire_l1_w0_n41_mux_dataout & wire_l1_w0_n40_mux_dataout
 & wire_l1_w0_n39_mux_dataout & wire_l1_w0_n38_mux_dataout & wire_l1_w0_n37_mux_dataout & wire_l1_w0_n36_mux_dataout & wire_l1_w0_n35_mux_dataout & wire_l1_w0_n34_mux_dataout & wire_l1_w0_n33_mux_dataout & wire_l1_w0_n32_mux_dataout & wire_l1_w0_n31_mux_dataout & wire_l1_w0_n30_mux_dataout & wire_l1_w0_n29_mux_dataout & wire_l1_w0_n28_mux_dataout & wire_l1_w0_n27_mux_dataout & wire_l1_w0_n26_mux_dataout & wire_l1_w0_n25_mux_dataout & wire_l1_w0_n24_mux_dataout & wire_l1_w0_n23_mux_dataout & wire_l1_w0_n22_mux_dataout & wire_l1_w0_n21_mux_dataout & wire_l1_w0_n20_mux_dataout & wire_l1_w0_n19_mux_dataout & wire_l1_w0_n18_mux_dataout & wire_l1_w0_n17_mux_dataout & wire_l1_w0_n16_mux_dataout & wire_l1_w0_n15_mux_dataout & wire_l1_w0_n14_mux_dataout & wire_l1_w0_n13_mux_dataout & wire_l1_w0_n12_mux_dataout & wire_l1_w0_n11_mux_dataout & wire_l1_w0_n10_mux_dataout & wire_l1_w0_n9_mux_dataout & wire_l1_w0_n8_mux_dataout & wire_l1_w0_n7_mux_dataout & wire_l1_w0_n6_mux_dataout & wire_l1_w0_n5_mux_dataout & wire_l1_w0_n4_mux_dataout & wire_l1_w0_n3_mux_dataout & wire_l1_w0_n2_mux_dataout & wire_l1_w0_n1_mux_dataout & wire_l1_w0_n0_mux_dataout & "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" & data);
	result <= result_wire_ext;
	result_wire_ext(0) <= ( wire_l8_w0_n0_mux_dataout);
	sel_wire <= ( sel(7) & "00000000" & sel(6) & "00000000" & sel(5) & "00000000" & sel(4) & "00000000" & sel(3) & "00000000" & sel(2) & "00000000" & sel(1) & "00000000" & sel(0));
	wire_l1_w0_n0_mux_dataout <= data_wire(1) WHEN sel_wire(0) = '1'  ELSE data_wire(0);
	wire_l1_w0_n100_mux_dataout <= data_wire(201) WHEN sel_wire(0) = '1'  ELSE data_wire(200);
	wire_l1_w0_n101_mux_dataout <= data_wire(203) WHEN sel_wire(0) = '1'  ELSE data_wire(202);
	wire_l1_w0_n102_mux_dataout <= data_wire(205) WHEN sel_wire(0) = '1'  ELSE data_wire(204);
	wire_l1_w0_n103_mux_dataout <= data_wire(207) WHEN sel_wire(0) = '1'  ELSE data_wire(206);
	wire_l1_w0_n104_mux_dataout <= data_wire(209) WHEN sel_wire(0) = '1'  ELSE data_wire(208);
	wire_l1_w0_n105_mux_dataout <= data_wire(211) WHEN sel_wire(0) = '1'  ELSE data_wire(210);
	wire_l1_w0_n106_mux_dataout <= data_wire(213) WHEN sel_wire(0) = '1'  ELSE data_wire(212);
	wire_l1_w0_n107_mux_dataout <= data_wire(215) WHEN sel_wire(0) = '1'  ELSE data_wire(214);
	wire_l1_w0_n108_mux_dataout <= data_wire(217) WHEN sel_wire(0) = '1'  ELSE data_wire(216);
	wire_l1_w0_n109_mux_dataout <= data_wire(219) WHEN sel_wire(0) = '1'  ELSE data_wire(218);
	wire_l1_w0_n10_mux_dataout <= data_wire(21) WHEN sel_wire(0) = '1'  ELSE data_wire(20);
	wire_l1_w0_n110_mux_dataout <= data_wire(221) WHEN sel_wire(0) = '1'  ELSE data_wire(220);
	wire_l1_w0_n111_mux_dataout <= data_wire(223) WHEN sel_wire(0) = '1'  ELSE data_wire(222);
	wire_l1_w0_n112_mux_dataout <= data_wire(225) WHEN sel_wire(0) = '1'  ELSE data_wire(224);
	wire_l1_w0_n113_mux_dataout <= data_wire(227) WHEN sel_wire(0) = '1'  ELSE data_wire(226);
	wire_l1_w0_n114_mux_dataout <= data_wire(229) WHEN sel_wire(0) = '1'  ELSE data_wire(228);
	wire_l1_w0_n115_mux_dataout <= data_wire(231) WHEN sel_wire(0) = '1'  ELSE data_wire(230);
	wire_l1_w0_n116_mux_dataout <= data_wire(233) WHEN sel_wire(0) = '1'  ELSE data_wire(232);
	wire_l1_w0_n117_mux_dataout <= data_wire(235) WHEN sel_wire(0) = '1'  ELSE data_wire(234);
	wire_l1_w0_n118_mux_dataout <= data_wire(237) WHEN sel_wire(0) = '1'  ELSE data_wire(236);
	wire_l1_w0_n119_mux_dataout <= data_wire(239) WHEN sel_wire(0) = '1'  ELSE data_wire(238);
	wire_l1_w0_n11_mux_dataout <= data_wire(23) WHEN sel_wire(0) = '1'  ELSE data_wire(22);
	wire_l1_w0_n120_mux_dataout <= data_wire(241) WHEN sel_wire(0) = '1'  ELSE data_wire(240);
	wire_l1_w0_n121_mux_dataout <= data_wire(243) WHEN sel_wire(0) = '1'  ELSE data_wire(242);
	wire_l1_w0_n122_mux_dataout <= data_wire(245) WHEN sel_wire(0) = '1'  ELSE data_wire(244);
	wire_l1_w0_n123_mux_dataout <= data_wire(247) WHEN sel_wire(0) = '1'  ELSE data_wire(246);
	wire_l1_w0_n124_mux_dataout <= data_wire(249) WHEN sel_wire(0) = '1'  ELSE data_wire(248);
	wire_l1_w0_n125_mux_dataout <= data_wire(251) WHEN sel_wire(0) = '1'  ELSE data_wire(250);
	wire_l1_w0_n126_mux_dataout <= data_wire(253) WHEN sel_wire(0) = '1'  ELSE data_wire(252);
	wire_l1_w0_n127_mux_dataout <= data_wire(255) WHEN sel_wire(0) = '1'  ELSE data_wire(254);
	wire_l1_w0_n12_mux_dataout <= data_wire(25) WHEN sel_wire(0) = '1'  ELSE data_wire(24);
	wire_l1_w0_n13_mux_dataout <= data_wire(27) WHEN sel_wire(0) = '1'  ELSE data_wire(26);
	wire_l1_w0_n14_mux_dataout <= data_wire(29) WHEN sel_wire(0) = '1'  ELSE data_wire(28);
	wire_l1_w0_n15_mux_dataout <= data_wire(31) WHEN sel_wire(0) = '1'  ELSE data_wire(30);
	wire_l1_w0_n16_mux_dataout <= data_wire(33) WHEN sel_wire(0) = '1'  ELSE data_wire(32);
	wire_l1_w0_n17_mux_dataout <= data_wire(35) WHEN sel_wire(0) = '1'  ELSE data_wire(34);
	wire_l1_w0_n18_mux_dataout <= data_wire(37) WHEN sel_wire(0) = '1'  ELSE data_wire(36);
	wire_l1_w0_n19_mux_dataout <= data_wire(39) WHEN sel_wire(0) = '1'  ELSE data_wire(38);
	wire_l1_w0_n1_mux_dataout <= data_wire(3) WHEN sel_wire(0) = '1'  ELSE data_wire(2);
	wire_l1_w0_n20_mux_dataout <= data_wire(41) WHEN sel_wire(0) = '1'  ELSE data_wire(40);
	wire_l1_w0_n21_mux_dataout <= data_wire(43) WHEN sel_wire(0) = '1'  ELSE data_wire(42);
	wire_l1_w0_n22_mux_dataout <= data_wire(45) WHEN sel_wire(0) = '1'  ELSE data_wire(44);
	wire_l1_w0_n23_mux_dataout <= data_wire(47) WHEN sel_wire(0) = '1'  ELSE data_wire(46);
	wire_l1_w0_n24_mux_dataout <= data_wire(49) WHEN sel_wire(0) = '1'  ELSE data_wire(48);
	wire_l1_w0_n25_mux_dataout <= data_wire(51) WHEN sel_wire(0) = '1'  ELSE data_wire(50);
	wire_l1_w0_n26_mux_dataout <= data_wire(53) WHEN sel_wire(0) = '1'  ELSE data_wire(52);
	wire_l1_w0_n27_mux_dataout <= data_wire(55) WHEN sel_wire(0) = '1'  ELSE data_wire(54);
	wire_l1_w0_n28_mux_dataout <= data_wire(57) WHEN sel_wire(0) = '1'  ELSE data_wire(56);
	wire_l1_w0_n29_mux_dataout <= data_wire(59) WHEN sel_wire(0) = '1'  ELSE data_wire(58);
	wire_l1_w0_n2_mux_dataout <= data_wire(5) WHEN sel_wire(0) = '1'  ELSE data_wire(4);
	wire_l1_w0_n30_mux_dataout <= data_wire(61) WHEN sel_wire(0) = '1'  ELSE data_wire(60);
	wire_l1_w0_n31_mux_dataout <= data_wire(63) WHEN sel_wire(0) = '1'  ELSE data_wire(62);
	wire_l1_w0_n32_mux_dataout <= data_wire(65) WHEN sel_wire(0) = '1'  ELSE data_wire(64);
	wire_l1_w0_n33_mux_dataout <= data_wire(67) WHEN sel_wire(0) = '1'  ELSE data_wire(66);
	wire_l1_w0_n34_mux_dataout <= data_wire(69) WHEN sel_wire(0) = '1'  ELSE data_wire(68);
	wire_l1_w0_n35_mux_dataout <= data_wire(71) WHEN sel_wire(0) = '1'  ELSE data_wire(70);
	wire_l1_w0_n36_mux_dataout <= data_wire(73) WHEN sel_wire(0) = '1'  ELSE data_wire(72);
	wire_l1_w0_n37_mux_dataout <= data_wire(75) WHEN sel_wire(0) = '1'  ELSE data_wire(74);
	wire_l1_w0_n38_mux_dataout <= data_wire(77) WHEN sel_wire(0) = '1'  ELSE data_wire(76);
	wire_l1_w0_n39_mux_dataout <= data_wire(79) WHEN sel_wire(0) = '1'  ELSE data_wire(78);
	wire_l1_w0_n3_mux_dataout <= data_wire(7) WHEN sel_wire(0) = '1'  ELSE data_wire(6);
	wire_l1_w0_n40_mux_dataout <= data_wire(81) WHEN sel_wire(0) = '1'  ELSE data_wire(80);
	wire_l1_w0_n41_mux_dataout <= data_wire(83) WHEN sel_wire(0) = '1'  ELSE data_wire(82);
	wire_l1_w0_n42_mux_dataout <= data_wire(85) WHEN sel_wire(0) = '1'  ELSE data_wire(84);
	wire_l1_w0_n43_mux_dataout <= data_wire(87) WHEN sel_wire(0) = '1'  ELSE data_wire(86);
	wire_l1_w0_n44_mux_dataout <= data_wire(89) WHEN sel_wire(0) = '1'  ELSE data_wire(88);
	wire_l1_w0_n45_mux_dataout <= data_wire(91) WHEN sel_wire(0) = '1'  ELSE data_wire(90);
	wire_l1_w0_n46_mux_dataout <= data_wire(93) WHEN sel_wire(0) = '1'  ELSE data_wire(92);
	wire_l1_w0_n47_mux_dataout <= data_wire(95) WHEN sel_wire(0) = '1'  ELSE data_wire(94);
	wire_l1_w0_n48_mux_dataout <= data_wire(97) WHEN sel_wire(0) = '1'  ELSE data_wire(96);
	wire_l1_w0_n49_mux_dataout <= data_wire(99) WHEN sel_wire(0) = '1'  ELSE data_wire(98);
	wire_l1_w0_n4_mux_dataout <= data_wire(9) WHEN sel_wire(0) = '1'  ELSE data_wire(8);
	wire_l1_w0_n50_mux_dataout <= data_wire(101) WHEN sel_wire(0) = '1'  ELSE data_wire(100);
	wire_l1_w0_n51_mux_dataout <= data_wire(103) WHEN sel_wire(0) = '1'  ELSE data_wire(102);
	wire_l1_w0_n52_mux_dataout <= data_wire(105) WHEN sel_wire(0) = '1'  ELSE data_wire(104);
	wire_l1_w0_n53_mux_dataout <= data_wire(107) WHEN sel_wire(0) = '1'  ELSE data_wire(106);
	wire_l1_w0_n54_mux_dataout <= data_wire(109) WHEN sel_wire(0) = '1'  ELSE data_wire(108);
	wire_l1_w0_n55_mux_dataout <= data_wire(111) WHEN sel_wire(0) = '1'  ELSE data_wire(110);
	wire_l1_w0_n56_mux_dataout <= data_wire(113) WHEN sel_wire(0) = '1'  ELSE data_wire(112);
	wire_l1_w0_n57_mux_dataout <= data_wire(115) WHEN sel_wire(0) = '1'  ELSE data_wire(114);
	wire_l1_w0_n58_mux_dataout <= data_wire(117) WHEN sel_wire(0) = '1'  ELSE data_wire(116);
	wire_l1_w0_n59_mux_dataout <= data_wire(119) WHEN sel_wire(0) = '1'  ELSE data_wire(118);
	wire_l1_w0_n5_mux_dataout <= data_wire(11) WHEN sel_wire(0) = '1'  ELSE data_wire(10);
	wire_l1_w0_n60_mux_dataout <= data_wire(121) WHEN sel_wire(0) = '1'  ELSE data_wire(120);
	wire_l1_w0_n61_mux_dataout <= data_wire(123) WHEN sel_wire(0) = '1'  ELSE data_wire(122);
	wire_l1_w0_n62_mux_dataout <= data_wire(125) WHEN sel_wire(0) = '1'  ELSE data_wire(124);
	wire_l1_w0_n63_mux_dataout <= data_wire(127) WHEN sel_wire(0) = '1'  ELSE data_wire(126);
	wire_l1_w0_n64_mux_dataout <= data_wire(129) WHEN sel_wire(0) = '1'  ELSE data_wire(128);
	wire_l1_w0_n65_mux_dataout <= data_wire(131) WHEN sel_wire(0) = '1'  ELSE data_wire(130);
	wire_l1_w0_n66_mux_dataout <= data_wire(133) WHEN sel_wire(0) = '1'  ELSE data_wire(132);
	wire_l1_w0_n67_mux_dataout <= data_wire(135) WHEN sel_wire(0) = '1'  ELSE data_wire(134);
	wire_l1_w0_n68_mux_dataout <= data_wire(137) WHEN sel_wire(0) = '1'  ELSE data_wire(136);
	wire_l1_w0_n69_mux_dataout <= data_wire(139) WHEN sel_wire(0) = '1'  ELSE data_wire(138);
	wire_l1_w0_n6_mux_dataout <= data_wire(13) WHEN sel_wire(0) = '1'  ELSE data_wire(12);
	wire_l1_w0_n70_mux_dataout <= data_wire(141) WHEN sel_wire(0) = '1'  ELSE data_wire(140);
	wire_l1_w0_n71_mux_dataout <= data_wire(143) WHEN sel_wire(0) = '1'  ELSE data_wire(142);
	wire_l1_w0_n72_mux_dataout <= data_wire(145) WHEN sel_wire(0) = '1'  ELSE data_wire(144);
	wire_l1_w0_n73_mux_dataout <= data_wire(147) WHEN sel_wire(0) = '1'  ELSE data_wire(146);
	wire_l1_w0_n74_mux_dataout <= data_wire(149) WHEN sel_wire(0) = '1'  ELSE data_wire(148);
	wire_l1_w0_n75_mux_dataout <= data_wire(151) WHEN sel_wire(0) = '1'  ELSE data_wire(150);
	wire_l1_w0_n76_mux_dataout <= data_wire(153) WHEN sel_wire(0) = '1'  ELSE data_wire(152);
	wire_l1_w0_n77_mux_dataout <= data_wire(155) WHEN sel_wire(0) = '1'  ELSE data_wire(154);
	wire_l1_w0_n78_mux_dataout <= data_wire(157) WHEN sel_wire(0) = '1'  ELSE data_wire(156);
	wire_l1_w0_n79_mux_dataout <= data_wire(159) WHEN sel_wire(0) = '1'  ELSE data_wire(158);
	wire_l1_w0_n7_mux_dataout <= data_wire(15) WHEN sel_wire(0) = '1'  ELSE data_wire(14);
	wire_l1_w0_n80_mux_dataout <= data_wire(161) WHEN sel_wire(0) = '1'  ELSE data_wire(160);
	wire_l1_w0_n81_mux_dataout <= data_wire(163) WHEN sel_wire(0) = '1'  ELSE data_wire(162);
	wire_l1_w0_n82_mux_dataout <= data_wire(165) WHEN sel_wire(0) = '1'  ELSE data_wire(164);
	wire_l1_w0_n83_mux_dataout <= data_wire(167) WHEN sel_wire(0) = '1'  ELSE data_wire(166);
	wire_l1_w0_n84_mux_dataout <= data_wire(169) WHEN sel_wire(0) = '1'  ELSE data_wire(168);
	wire_l1_w0_n85_mux_dataout <= data_wire(171) WHEN sel_wire(0) = '1'  ELSE data_wire(170);
	wire_l1_w0_n86_mux_dataout <= data_wire(173) WHEN sel_wire(0) = '1'  ELSE data_wire(172);
	wire_l1_w0_n87_mux_dataout <= data_wire(175) WHEN sel_wire(0) = '1'  ELSE data_wire(174);
	wire_l1_w0_n88_mux_dataout <= data_wire(177) WHEN sel_wire(0) = '1'  ELSE data_wire(176);
	wire_l1_w0_n89_mux_dataout <= data_wire(179) WHEN sel_wire(0) = '1'  ELSE data_wire(178);
	wire_l1_w0_n8_mux_dataout <= data_wire(17) WHEN sel_wire(0) = '1'  ELSE data_wire(16);
	wire_l1_w0_n90_mux_dataout <= data_wire(181) WHEN sel_wire(0) = '1'  ELSE data_wire(180);
	wire_l1_w0_n91_mux_dataout <= data_wire(183) WHEN sel_wire(0) = '1'  ELSE data_wire(182);
	wire_l1_w0_n92_mux_dataout <= data_wire(185) WHEN sel_wire(0) = '1'  ELSE data_wire(184);
	wire_l1_w0_n93_mux_dataout <= data_wire(187) WHEN sel_wire(0) = '1'  ELSE data_wire(186);
	wire_l1_w0_n94_mux_dataout <= data_wire(189) WHEN sel_wire(0) = '1'  ELSE data_wire(188);
	wire_l1_w0_n95_mux_dataout <= data_wire(191) WHEN sel_wire(0) = '1'  ELSE data_wire(190);
	wire_l1_w0_n96_mux_dataout <= data_wire(193) WHEN sel_wire(0) = '1'  ELSE data_wire(192);
	wire_l1_w0_n97_mux_dataout <= data_wire(195) WHEN sel_wire(0) = '1'  ELSE data_wire(194);
	wire_l1_w0_n98_mux_dataout <= data_wire(197) WHEN sel_wire(0) = '1'  ELSE data_wire(196);
	wire_l1_w0_n99_mux_dataout <= data_wire(199) WHEN sel_wire(0) = '1'  ELSE data_wire(198);
	wire_l1_w0_n9_mux_dataout <= data_wire(19) WHEN sel_wire(0) = '1'  ELSE data_wire(18);
	wire_l2_w0_n0_mux_dataout <= data_wire(257) WHEN sel_wire(9) = '1'  ELSE data_wire(256);
	wire_l2_w0_n10_mux_dataout <= data_wire(277) WHEN sel_wire(9) = '1'  ELSE data_wire(276);
	wire_l2_w0_n11_mux_dataout <= data_wire(279) WHEN sel_wire(9) = '1'  ELSE data_wire(278);
	wire_l2_w0_n12_mux_dataout <= data_wire(281) WHEN sel_wire(9) = '1'  ELSE data_wire(280);
	wire_l2_w0_n13_mux_dataout <= data_wire(283) WHEN sel_wire(9) = '1'  ELSE data_wire(282);
	wire_l2_w0_n14_mux_dataout <= data_wire(285) WHEN sel_wire(9) = '1'  ELSE data_wire(284);
	wire_l2_w0_n15_mux_dataout <= data_wire(287) WHEN sel_wire(9) = '1'  ELSE data_wire(286);
	wire_l2_w0_n16_mux_dataout <= data_wire(289) WHEN sel_wire(9) = '1'  ELSE data_wire(288);
	wire_l2_w0_n17_mux_dataout <= data_wire(291) WHEN sel_wire(9) = '1'  ELSE data_wire(290);
	wire_l2_w0_n18_mux_dataout <= data_wire(293) WHEN sel_wire(9) = '1'  ELSE data_wire(292);
	wire_l2_w0_n19_mux_dataout <= data_wire(295) WHEN sel_wire(9) = '1'  ELSE data_wire(294);
	wire_l2_w0_n1_mux_dataout <= data_wire(259) WHEN sel_wire(9) = '1'  ELSE data_wire(258);
	wire_l2_w0_n20_mux_dataout <= data_wire(297) WHEN sel_wire(9) = '1'  ELSE data_wire(296);
	wire_l2_w0_n21_mux_dataout <= data_wire(299) WHEN sel_wire(9) = '1'  ELSE data_wire(298);
	wire_l2_w0_n22_mux_dataout <= data_wire(301) WHEN sel_wire(9) = '1'  ELSE data_wire(300);
	wire_l2_w0_n23_mux_dataout <= data_wire(303) WHEN sel_wire(9) = '1'  ELSE data_wire(302);
	wire_l2_w0_n24_mux_dataout <= data_wire(305) WHEN sel_wire(9) = '1'  ELSE data_wire(304);
	wire_l2_w0_n25_mux_dataout <= data_wire(307) WHEN sel_wire(9) = '1'  ELSE data_wire(306);
	wire_l2_w0_n26_mux_dataout <= data_wire(309) WHEN sel_wire(9) = '1'  ELSE data_wire(308);
	wire_l2_w0_n27_mux_dataout <= data_wire(311) WHEN sel_wire(9) = '1'  ELSE data_wire(310);
	wire_l2_w0_n28_mux_dataout <= data_wire(313) WHEN sel_wire(9) = '1'  ELSE data_wire(312);
	wire_l2_w0_n29_mux_dataout <= data_wire(315) WHEN sel_wire(9) = '1'  ELSE data_wire(314);
	wire_l2_w0_n2_mux_dataout <= data_wire(261) WHEN sel_wire(9) = '1'  ELSE data_wire(260);
	wire_l2_w0_n30_mux_dataout <= data_wire(317) WHEN sel_wire(9) = '1'  ELSE data_wire(316);
	wire_l2_w0_n31_mux_dataout <= data_wire(319) WHEN sel_wire(9) = '1'  ELSE data_wire(318);
	wire_l2_w0_n32_mux_dataout <= data_wire(321) WHEN sel_wire(9) = '1'  ELSE data_wire(320);
	wire_l2_w0_n33_mux_dataout <= data_wire(323) WHEN sel_wire(9) = '1'  ELSE data_wire(322);
	wire_l2_w0_n34_mux_dataout <= data_wire(325) WHEN sel_wire(9) = '1'  ELSE data_wire(324);
	wire_l2_w0_n35_mux_dataout <= data_wire(327) WHEN sel_wire(9) = '1'  ELSE data_wire(326);
	wire_l2_w0_n36_mux_dataout <= data_wire(329) WHEN sel_wire(9) = '1'  ELSE data_wire(328);
	wire_l2_w0_n37_mux_dataout <= data_wire(331) WHEN sel_wire(9) = '1'  ELSE data_wire(330);
	wire_l2_w0_n38_mux_dataout <= data_wire(333) WHEN sel_wire(9) = '1'  ELSE data_wire(332);
	wire_l2_w0_n39_mux_dataout <= data_wire(335) WHEN sel_wire(9) = '1'  ELSE data_wire(334);
	wire_l2_w0_n3_mux_dataout <= data_wire(263) WHEN sel_wire(9) = '1'  ELSE data_wire(262);
	wire_l2_w0_n40_mux_dataout <= data_wire(337) WHEN sel_wire(9) = '1'  ELSE data_wire(336);
	wire_l2_w0_n41_mux_dataout <= data_wire(339) WHEN sel_wire(9) = '1'  ELSE data_wire(338);
	wire_l2_w0_n42_mux_dataout <= data_wire(341) WHEN sel_wire(9) = '1'  ELSE data_wire(340);
	wire_l2_w0_n43_mux_dataout <= data_wire(343) WHEN sel_wire(9) = '1'  ELSE data_wire(342);
	wire_l2_w0_n44_mux_dataout <= data_wire(345) WHEN sel_wire(9) = '1'  ELSE data_wire(344);
	wire_l2_w0_n45_mux_dataout <= data_wire(347) WHEN sel_wire(9) = '1'  ELSE data_wire(346);
	wire_l2_w0_n46_mux_dataout <= data_wire(349) WHEN sel_wire(9) = '1'  ELSE data_wire(348);
	wire_l2_w0_n47_mux_dataout <= data_wire(351) WHEN sel_wire(9) = '1'  ELSE data_wire(350);
	wire_l2_w0_n48_mux_dataout <= data_wire(353) WHEN sel_wire(9) = '1'  ELSE data_wire(352);
	wire_l2_w0_n49_mux_dataout <= data_wire(355) WHEN sel_wire(9) = '1'  ELSE data_wire(354);
	wire_l2_w0_n4_mux_dataout <= data_wire(265) WHEN sel_wire(9) = '1'  ELSE data_wire(264);
	wire_l2_w0_n50_mux_dataout <= data_wire(357) WHEN sel_wire(9) = '1'  ELSE data_wire(356);
	wire_l2_w0_n51_mux_dataout <= data_wire(359) WHEN sel_wire(9) = '1'  ELSE data_wire(358);
	wire_l2_w0_n52_mux_dataout <= data_wire(361) WHEN sel_wire(9) = '1'  ELSE data_wire(360);
	wire_l2_w0_n53_mux_dataout <= data_wire(363) WHEN sel_wire(9) = '1'  ELSE data_wire(362);
	wire_l2_w0_n54_mux_dataout <= data_wire(365) WHEN sel_wire(9) = '1'  ELSE data_wire(364);
	wire_l2_w0_n55_mux_dataout <= data_wire(367) WHEN sel_wire(9) = '1'  ELSE data_wire(366);
	wire_l2_w0_n56_mux_dataout <= data_wire(369) WHEN sel_wire(9) = '1'  ELSE data_wire(368);
	wire_l2_w0_n57_mux_dataout <= data_wire(371) WHEN sel_wire(9) = '1'  ELSE data_wire(370);
	wire_l2_w0_n58_mux_dataout <= data_wire(373) WHEN sel_wire(9) = '1'  ELSE data_wire(372);
	wire_l2_w0_n59_mux_dataout <= data_wire(375) WHEN sel_wire(9) = '1'  ELSE data_wire(374);
	wire_l2_w0_n5_mux_dataout <= data_wire(267) WHEN sel_wire(9) = '1'  ELSE data_wire(266);
	wire_l2_w0_n60_mux_dataout <= data_wire(377) WHEN sel_wire(9) = '1'  ELSE data_wire(376);
	wire_l2_w0_n61_mux_dataout <= data_wire(379) WHEN sel_wire(9) = '1'  ELSE data_wire(378);
	wire_l2_w0_n62_mux_dataout <= data_wire(381) WHEN sel_wire(9) = '1'  ELSE data_wire(380);
	wire_l2_w0_n63_mux_dataout <= data_wire(383) WHEN sel_wire(9) = '1'  ELSE data_wire(382);
	wire_l2_w0_n6_mux_dataout <= data_wire(269) WHEN sel_wire(9) = '1'  ELSE data_wire(268);
	wire_l2_w0_n7_mux_dataout <= data_wire(271) WHEN sel_wire(9) = '1'  ELSE data_wire(270);
	wire_l2_w0_n8_mux_dataout <= data_wire(273) WHEN sel_wire(9) = '1'  ELSE data_wire(272);
	wire_l2_w0_n9_mux_dataout <= data_wire(275) WHEN sel_wire(9) = '1'  ELSE data_wire(274);
	wire_l3_w0_n0_mux_dataout <= data_wire(385) WHEN sel_wire(18) = '1'  ELSE data_wire(384);
	wire_l3_w0_n10_mux_dataout <= data_wire(405) WHEN sel_wire(18) = '1'  ELSE data_wire(404);
	wire_l3_w0_n11_mux_dataout <= data_wire(407) WHEN sel_wire(18) = '1'  ELSE data_wire(406);
	wire_l3_w0_n12_mux_dataout <= data_wire(409) WHEN sel_wire(18) = '1'  ELSE data_wire(408);
	wire_l3_w0_n13_mux_dataout <= data_wire(411) WHEN sel_wire(18) = '1'  ELSE data_wire(410);
	wire_l3_w0_n14_mux_dataout <= data_wire(413) WHEN sel_wire(18) = '1'  ELSE data_wire(412);
	wire_l3_w0_n15_mux_dataout <= data_wire(415) WHEN sel_wire(18) = '1'  ELSE data_wire(414);
	wire_l3_w0_n16_mux_dataout <= data_wire(417) WHEN sel_wire(18) = '1'  ELSE data_wire(416);
	wire_l3_w0_n17_mux_dataout <= data_wire(419) WHEN sel_wire(18) = '1'  ELSE data_wire(418);
	wire_l3_w0_n18_mux_dataout <= data_wire(421) WHEN sel_wire(18) = '1'  ELSE data_wire(420);
	wire_l3_w0_n19_mux_dataout <= data_wire(423) WHEN sel_wire(18) = '1'  ELSE data_wire(422);
	wire_l3_w0_n1_mux_dataout <= data_wire(387) WHEN sel_wire(18) = '1'  ELSE data_wire(386);
	wire_l3_w0_n20_mux_dataout <= data_wire(425) WHEN sel_wire(18) = '1'  ELSE data_wire(424);
	wire_l3_w0_n21_mux_dataout <= data_wire(427) WHEN sel_wire(18) = '1'  ELSE data_wire(426);
	wire_l3_w0_n22_mux_dataout <= data_wire(429) WHEN sel_wire(18) = '1'  ELSE data_wire(428);
	wire_l3_w0_n23_mux_dataout <= data_wire(431) WHEN sel_wire(18) = '1'  ELSE data_wire(430);
	wire_l3_w0_n24_mux_dataout <= data_wire(433) WHEN sel_wire(18) = '1'  ELSE data_wire(432);
	wire_l3_w0_n25_mux_dataout <= data_wire(435) WHEN sel_wire(18) = '1'  ELSE data_wire(434);
	wire_l3_w0_n26_mux_dataout <= data_wire(437) WHEN sel_wire(18) = '1'  ELSE data_wire(436);
	wire_l3_w0_n27_mux_dataout <= data_wire(439) WHEN sel_wire(18) = '1'  ELSE data_wire(438);
	wire_l3_w0_n28_mux_dataout <= data_wire(441) WHEN sel_wire(18) = '1'  ELSE data_wire(440);
	wire_l3_w0_n29_mux_dataout <= data_wire(443) WHEN sel_wire(18) = '1'  ELSE data_wire(442);
	wire_l3_w0_n2_mux_dataout <= data_wire(389) WHEN sel_wire(18) = '1'  ELSE data_wire(388);
	wire_l3_w0_n30_mux_dataout <= data_wire(445) WHEN sel_wire(18) = '1'  ELSE data_wire(444);
	wire_l3_w0_n31_mux_dataout <= data_wire(447) WHEN sel_wire(18) = '1'  ELSE data_wire(446);
	wire_l3_w0_n3_mux_dataout <= data_wire(391) WHEN sel_wire(18) = '1'  ELSE data_wire(390);
	wire_l3_w0_n4_mux_dataout <= data_wire(393) WHEN sel_wire(18) = '1'  ELSE data_wire(392);
	wire_l3_w0_n5_mux_dataout <= data_wire(395) WHEN sel_wire(18) = '1'  ELSE data_wire(394);
	wire_l3_w0_n6_mux_dataout <= data_wire(397) WHEN sel_wire(18) = '1'  ELSE data_wire(396);
	wire_l3_w0_n7_mux_dataout <= data_wire(399) WHEN sel_wire(18) = '1'  ELSE data_wire(398);
	wire_l3_w0_n8_mux_dataout <= data_wire(401) WHEN sel_wire(18) = '1'  ELSE data_wire(400);
	wire_l3_w0_n9_mux_dataout <= data_wire(403) WHEN sel_wire(18) = '1'  ELSE data_wire(402);
	wire_l4_w0_n0_mux_dataout <= data_wire(449) WHEN sel_wire(27) = '1'  ELSE data_wire(448);
	wire_l4_w0_n10_mux_dataout <= data_wire(469) WHEN sel_wire(27) = '1'  ELSE data_wire(468);
	wire_l4_w0_n11_mux_dataout <= data_wire(471) WHEN sel_wire(27) = '1'  ELSE data_wire(470);
	wire_l4_w0_n12_mux_dataout <= data_wire(473) WHEN sel_wire(27) = '1'  ELSE data_wire(472);
	wire_l4_w0_n13_mux_dataout <= data_wire(475) WHEN sel_wire(27) = '1'  ELSE data_wire(474);
	wire_l4_w0_n14_mux_dataout <= data_wire(477) WHEN sel_wire(27) = '1'  ELSE data_wire(476);
	wire_l4_w0_n15_mux_dataout <= data_wire(479) WHEN sel_wire(27) = '1'  ELSE data_wire(478);
	wire_l4_w0_n1_mux_dataout <= data_wire(451) WHEN sel_wire(27) = '1'  ELSE data_wire(450);
	wire_l4_w0_n2_mux_dataout <= data_wire(453) WHEN sel_wire(27) = '1'  ELSE data_wire(452);
	wire_l4_w0_n3_mux_dataout <= data_wire(455) WHEN sel_wire(27) = '1'  ELSE data_wire(454);
	wire_l4_w0_n4_mux_dataout <= data_wire(457) WHEN sel_wire(27) = '1'  ELSE data_wire(456);
	wire_l4_w0_n5_mux_dataout <= data_wire(459) WHEN sel_wire(27) = '1'  ELSE data_wire(458);
	wire_l4_w0_n6_mux_dataout <= data_wire(461) WHEN sel_wire(27) = '1'  ELSE data_wire(460);
	wire_l4_w0_n7_mux_dataout <= data_wire(463) WHEN sel_wire(27) = '1'  ELSE data_wire(462);
	wire_l4_w0_n8_mux_dataout <= data_wire(465) WHEN sel_wire(27) = '1'  ELSE data_wire(464);
	wire_l4_w0_n9_mux_dataout <= data_wire(467) WHEN sel_wire(27) = '1'  ELSE data_wire(466);
	wire_l5_w0_n0_mux_dataout <= data_wire(481) WHEN sel_wire(36) = '1'  ELSE data_wire(480);
	wire_l5_w0_n1_mux_dataout <= data_wire(483) WHEN sel_wire(36) = '1'  ELSE data_wire(482);
	wire_l5_w0_n2_mux_dataout <= data_wire(485) WHEN sel_wire(36) = '1'  ELSE data_wire(484);
	wire_l5_w0_n3_mux_dataout <= data_wire(487) WHEN sel_wire(36) = '1'  ELSE data_wire(486);
	wire_l5_w0_n4_mux_dataout <= data_wire(489) WHEN sel_wire(36) = '1'  ELSE data_wire(488);
	wire_l5_w0_n5_mux_dataout <= data_wire(491) WHEN sel_wire(36) = '1'  ELSE data_wire(490);
	wire_l5_w0_n6_mux_dataout <= data_wire(493) WHEN sel_wire(36) = '1'  ELSE data_wire(492);
	wire_l5_w0_n7_mux_dataout <= data_wire(495) WHEN sel_wire(36) = '1'  ELSE data_wire(494);
	wire_l6_w0_n0_mux_dataout <= data_wire(497) WHEN sel_wire(45) = '1'  ELSE data_wire(496);
	wire_l6_w0_n1_mux_dataout <= data_wire(499) WHEN sel_wire(45) = '1'  ELSE data_wire(498);
	wire_l6_w0_n2_mux_dataout <= data_wire(501) WHEN sel_wire(45) = '1'  ELSE data_wire(500);
	wire_l6_w0_n3_mux_dataout <= data_wire(503) WHEN sel_wire(45) = '1'  ELSE data_wire(502);
	wire_l7_w0_n0_mux_dataout <= data_wire(505) WHEN sel_wire(54) = '1'  ELSE data_wire(504);
	wire_l7_w0_n1_mux_dataout <= data_wire(507) WHEN sel_wire(54) = '1'  ELSE data_wire(506);
	wire_l8_w0_n0_mux_dataout <= data_wire(509) WHEN sel_wire(63) = '1'  ELSE data_wire(508);

 END RTL; --reconfig_side_mux_i9a


--lpm_mux CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix IV" LPM_SIZE=36 LPM_WIDTH=1 LPM_WIDTHS=6 data result sel
--VERSION_BEGIN 13.0 cbx_lpm_mux 2013:06:12:18:03:33:SJ cbx_mgl 2013:06:12:18:33:59:SJ  VERSION_END

--synthesis_resources = lut 21 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  reconfig_side_mux_08a IS 
	 PORT 
	 ( 
		 data	:	IN  STD_LOGIC_VECTOR (35 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (0 DOWNTO 0);
		 sel	:	IN  STD_LOGIC_VECTOR (5 DOWNTO 0) := (OTHERS => '0')
	 ); 
 END reconfig_side_mux_08a;

 ARCHITECTURE RTL OF reconfig_side_mux_08a IS

	 SIGNAL	wire_l1_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n10_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n11_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n12_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n13_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n14_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n15_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n16_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n17_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n18_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n19_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n20_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n21_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n22_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n23_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n24_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n25_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n26_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n27_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n28_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n29_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n30_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n31_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n4_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n5_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n6_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n7_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n8_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l1_w0_n9_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n10_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n11_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n12_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n13_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n14_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n15_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n4_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n5_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n6_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n7_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n8_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l2_w0_n9_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n4_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n5_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n6_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l3_w0_n7_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n2_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l4_w0_n3_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l5_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l5_w0_n1_mux_dataout	:	STD_LOGIC;
	 SIGNAL	wire_l6_w0_n0_mux_dataout	:	STD_LOGIC;
	 SIGNAL  data_wire :	STD_LOGIC_VECTOR (125 DOWNTO 0);
	 SIGNAL  result_wire_ext :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  sel_wire :	STD_LOGIC_VECTOR (35 DOWNTO 0);
 BEGIN

	data_wire <= ( wire_l5_w0_n1_mux_dataout & wire_l5_w0_n0_mux_dataout & wire_l4_w0_n3_mux_dataout & wire_l4_w0_n2_mux_dataout & wire_l4_w0_n1_mux_dataout & wire_l4_w0_n0_mux_dataout & wire_l3_w0_n7_mux_dataout & wire_l3_w0_n6_mux_dataout & wire_l3_w0_n5_mux_dataout & wire_l3_w0_n4_mux_dataout & wire_l3_w0_n3_mux_dataout & wire_l3_w0_n2_mux_dataout & wire_l3_w0_n1_mux_dataout & wire_l3_w0_n0_mux_dataout & wire_l2_w0_n15_mux_dataout & wire_l2_w0_n14_mux_dataout & wire_l2_w0_n13_mux_dataout & wire_l2_w0_n12_mux_dataout & wire_l2_w0_n11_mux_dataout & wire_l2_w0_n10_mux_dataout & wire_l2_w0_n9_mux_dataout & wire_l2_w0_n8_mux_dataout & wire_l2_w0_n7_mux_dataout & wire_l2_w0_n6_mux_dataout & wire_l2_w0_n5_mux_dataout & wire_l2_w0_n4_mux_dataout & wire_l2_w0_n3_mux_dataout & wire_l2_w0_n2_mux_dataout & wire_l2_w0_n1_mux_dataout & wire_l2_w0_n0_mux_dataout & wire_l1_w0_n31_mux_dataout & wire_l1_w0_n30_mux_dataout & wire_l1_w0_n29_mux_dataout & wire_l1_w0_n28_mux_dataout & wire_l1_w0_n27_mux_dataout & wire_l1_w0_n26_mux_dataout & wire_l1_w0_n25_mux_dataout & wire_l1_w0_n24_mux_dataout & wire_l1_w0_n23_mux_dataout & wire_l1_w0_n22_mux_dataout & wire_l1_w0_n21_mux_dataout & wire_l1_w0_n20_mux_dataout & wire_l1_w0_n19_mux_dataout & wire_l1_w0_n18_mux_dataout & wire_l1_w0_n17_mux_dataout & wire_l1_w0_n16_mux_dataout & wire_l1_w0_n15_mux_dataout & wire_l1_w0_n14_mux_dataout & wire_l1_w0_n13_mux_dataout & wire_l1_w0_n12_mux_dataout & wire_l1_w0_n11_mux_dataout & wire_l1_w0_n10_mux_dataout & wire_l1_w0_n9_mux_dataout & wire_l1_w0_n8_mux_dataout & wire_l1_w0_n7_mux_dataout & wire_l1_w0_n6_mux_dataout & wire_l1_w0_n5_mux_dataout & wire_l1_w0_n4_mux_dataout & wire_l1_w0_n3_mux_dataout & wire_l1_w0_n2_mux_dataout & wire_l1_w0_n1_mux_dataout & wire_l1_w0_n0_mux_dataout & "0000000000000000000000000000" & data);
	result <= result_wire_ext;
	result_wire_ext(0) <= ( wire_l6_w0_n0_mux_dataout);
	sel_wire <= ( sel(5) & "000000" & sel(4) & "000000" & sel(3) & "000000" & sel(2) & "000000" & sel(1) & "000000" & sel(0));
	wire_l1_w0_n0_mux_dataout <= data_wire(1) WHEN sel_wire(0) = '1'  ELSE data_wire(0);
	wire_l1_w0_n10_mux_dataout <= data_wire(21) WHEN sel_wire(0) = '1'  ELSE data_wire(20);
	wire_l1_w0_n11_mux_dataout <= data_wire(23) WHEN sel_wire(0) = '1'  ELSE data_wire(22);
	wire_l1_w0_n12_mux_dataout <= data_wire(25) WHEN sel_wire(0) = '1'  ELSE data_wire(24);
	wire_l1_w0_n13_mux_dataout <= data_wire(27) WHEN sel_wire(0) = '1'  ELSE data_wire(26);
	wire_l1_w0_n14_mux_dataout <= data_wire(29) WHEN sel_wire(0) = '1'  ELSE data_wire(28);
	wire_l1_w0_n15_mux_dataout <= data_wire(31) WHEN sel_wire(0) = '1'  ELSE data_wire(30);
	wire_l1_w0_n16_mux_dataout <= data_wire(33) WHEN sel_wire(0) = '1'  ELSE data_wire(32);
	wire_l1_w0_n17_mux_dataout <= data_wire(35) WHEN sel_wire(0) = '1'  ELSE data_wire(34);
	wire_l1_w0_n18_mux_dataout <= data_wire(37) WHEN sel_wire(0) = '1'  ELSE data_wire(36);
	wire_l1_w0_n19_mux_dataout <= data_wire(39) WHEN sel_wire(0) = '1'  ELSE data_wire(38);
	wire_l1_w0_n1_mux_dataout <= data_wire(3) WHEN sel_wire(0) = '1'  ELSE data_wire(2);
	wire_l1_w0_n20_mux_dataout <= data_wire(41) WHEN sel_wire(0) = '1'  ELSE data_wire(40);
	wire_l1_w0_n21_mux_dataout <= data_wire(43) WHEN sel_wire(0) = '1'  ELSE data_wire(42);
	wire_l1_w0_n22_mux_dataout <= data_wire(45) WHEN sel_wire(0) = '1'  ELSE data_wire(44);
	wire_l1_w0_n23_mux_dataout <= data_wire(47) WHEN sel_wire(0) = '1'  ELSE data_wire(46);
	wire_l1_w0_n24_mux_dataout <= data_wire(49) WHEN sel_wire(0) = '1'  ELSE data_wire(48);
	wire_l1_w0_n25_mux_dataout <= data_wire(51) WHEN sel_wire(0) = '1'  ELSE data_wire(50);
	wire_l1_w0_n26_mux_dataout <= data_wire(53) WHEN sel_wire(0) = '1'  ELSE data_wire(52);
	wire_l1_w0_n27_mux_dataout <= data_wire(55) WHEN sel_wire(0) = '1'  ELSE data_wire(54);
	wire_l1_w0_n28_mux_dataout <= data_wire(57) WHEN sel_wire(0) = '1'  ELSE data_wire(56);
	wire_l1_w0_n29_mux_dataout <= data_wire(59) WHEN sel_wire(0) = '1'  ELSE data_wire(58);
	wire_l1_w0_n2_mux_dataout <= data_wire(5) WHEN sel_wire(0) = '1'  ELSE data_wire(4);
	wire_l1_w0_n30_mux_dataout <= data_wire(61) WHEN sel_wire(0) = '1'  ELSE data_wire(60);
	wire_l1_w0_n31_mux_dataout <= data_wire(63) WHEN sel_wire(0) = '1'  ELSE data_wire(62);
	wire_l1_w0_n3_mux_dataout <= data_wire(7) WHEN sel_wire(0) = '1'  ELSE data_wire(6);
	wire_l1_w0_n4_mux_dataout <= data_wire(9) WHEN sel_wire(0) = '1'  ELSE data_wire(8);
	wire_l1_w0_n5_mux_dataout <= data_wire(11) WHEN sel_wire(0) = '1'  ELSE data_wire(10);
	wire_l1_w0_n6_mux_dataout <= data_wire(13) WHEN sel_wire(0) = '1'  ELSE data_wire(12);
	wire_l1_w0_n7_mux_dataout <= data_wire(15) WHEN sel_wire(0) = '1'  ELSE data_wire(14);
	wire_l1_w0_n8_mux_dataout <= data_wire(17) WHEN sel_wire(0) = '1'  ELSE data_wire(16);
	wire_l1_w0_n9_mux_dataout <= data_wire(19) WHEN sel_wire(0) = '1'  ELSE data_wire(18);
	wire_l2_w0_n0_mux_dataout <= data_wire(65) WHEN sel_wire(7) = '1'  ELSE data_wire(64);
	wire_l2_w0_n10_mux_dataout <= data_wire(85) WHEN sel_wire(7) = '1'  ELSE data_wire(84);
	wire_l2_w0_n11_mux_dataout <= data_wire(87) WHEN sel_wire(7) = '1'  ELSE data_wire(86);
	wire_l2_w0_n12_mux_dataout <= data_wire(89) WHEN sel_wire(7) = '1'  ELSE data_wire(88);
	wire_l2_w0_n13_mux_dataout <= data_wire(91) WHEN sel_wire(7) = '1'  ELSE data_wire(90);
	wire_l2_w0_n14_mux_dataout <= data_wire(93) WHEN sel_wire(7) = '1'  ELSE data_wire(92);
	wire_l2_w0_n15_mux_dataout <= data_wire(95) WHEN sel_wire(7) = '1'  ELSE data_wire(94);
	wire_l2_w0_n1_mux_dataout <= data_wire(67) WHEN sel_wire(7) = '1'  ELSE data_wire(66);
	wire_l2_w0_n2_mux_dataout <= data_wire(69) WHEN sel_wire(7) = '1'  ELSE data_wire(68);
	wire_l2_w0_n3_mux_dataout <= data_wire(71) WHEN sel_wire(7) = '1'  ELSE data_wire(70);
	wire_l2_w0_n4_mux_dataout <= data_wire(73) WHEN sel_wire(7) = '1'  ELSE data_wire(72);
	wire_l2_w0_n5_mux_dataout <= data_wire(75) WHEN sel_wire(7) = '1'  ELSE data_wire(74);
	wire_l2_w0_n6_mux_dataout <= data_wire(77) WHEN sel_wire(7) = '1'  ELSE data_wire(76);
	wire_l2_w0_n7_mux_dataout <= data_wire(79) WHEN sel_wire(7) = '1'  ELSE data_wire(78);
	wire_l2_w0_n8_mux_dataout <= data_wire(81) WHEN sel_wire(7) = '1'  ELSE data_wire(80);
	wire_l2_w0_n9_mux_dataout <= data_wire(83) WHEN sel_wire(7) = '1'  ELSE data_wire(82);
	wire_l3_w0_n0_mux_dataout <= data_wire(97) WHEN sel_wire(14) = '1'  ELSE data_wire(96);
	wire_l3_w0_n1_mux_dataout <= data_wire(99) WHEN sel_wire(14) = '1'  ELSE data_wire(98);
	wire_l3_w0_n2_mux_dataout <= data_wire(101) WHEN sel_wire(14) = '1'  ELSE data_wire(100);
	wire_l3_w0_n3_mux_dataout <= data_wire(103) WHEN sel_wire(14) = '1'  ELSE data_wire(102);
	wire_l3_w0_n4_mux_dataout <= data_wire(105) WHEN sel_wire(14) = '1'  ELSE data_wire(104);
	wire_l3_w0_n5_mux_dataout <= data_wire(107) WHEN sel_wire(14) = '1'  ELSE data_wire(106);
	wire_l3_w0_n6_mux_dataout <= data_wire(109) WHEN sel_wire(14) = '1'  ELSE data_wire(108);
	wire_l3_w0_n7_mux_dataout <= data_wire(111) WHEN sel_wire(14) = '1'  ELSE data_wire(110);
	wire_l4_w0_n0_mux_dataout <= data_wire(113) WHEN sel_wire(21) = '1'  ELSE data_wire(112);
	wire_l4_w0_n1_mux_dataout <= data_wire(115) WHEN sel_wire(21) = '1'  ELSE data_wire(114);
	wire_l4_w0_n2_mux_dataout <= data_wire(117) WHEN sel_wire(21) = '1'  ELSE data_wire(116);
	wire_l4_w0_n3_mux_dataout <= data_wire(119) WHEN sel_wire(21) = '1'  ELSE data_wire(118);
	wire_l5_w0_n0_mux_dataout <= data_wire(121) WHEN sel_wire(28) = '1'  ELSE data_wire(120);
	wire_l5_w0_n1_mux_dataout <= data_wire(123) WHEN sel_wire(28) = '1'  ELSE data_wire(122);
	wire_l6_w0_n0_mux_dataout <= data_wire(125) WHEN sel_wire(35) = '1'  ELSE data_wire(124);

 END RTL; --reconfig_side_mux_08a

 LIBRARY altera_mf;
 USE altera_mf.all;

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = alt_cal 1 alt_dfe 1 alt_eyemon 1 lpm_add_sub 4 lpm_compare 8 lpm_counter 5 lpm_decode 3 lut 153 reg 153 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  reconfig_side_alt2gxb_reconfig_4og2 IS 
	 PORT 
	 ( 
		 busy	:	OUT  STD_LOGIC;
		 ctrl_address	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
		 ctrl_read	:	IN  STD_LOGIC := '0';
		 ctrl_readdata	:	OUT  STD_LOGIC_VECTOR (15 DOWNTO 0);
		 ctrl_waitrequest	:	OUT  STD_LOGIC;
		 ctrl_write	:	IN  STD_LOGIC := '0';
		 ctrl_writedata	:	IN  STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
		 data_valid	:	OUT  STD_LOGIC;
		 error	:	OUT  STD_LOGIC;
		 logical_channel_address	:	IN  STD_LOGIC_VECTOR (7 DOWNTO 0) := (OTHERS => '0');
		 read	:	IN  STD_LOGIC := '0';
		 reconfig_clk	:	IN  STD_LOGIC;
		 reconfig_fromgxb	:	IN  STD_LOGIC_VECTOR (611 DOWNTO 0);
		 reconfig_mode_sel	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
		 reconfig_togxb	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 rx_eqctrl	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
		 rx_eqctrl_out	:	OUT  STD_LOGIC_VECTOR (3 DOWNTO 0);
		 rx_eqdcgain	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0');
		 rx_eqdcgain_out	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 tx_preemp_0t	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0) := (OTHERS => '0');
		 tx_preemp_0t_out	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 tx_preemp_1t	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0) := (OTHERS => '0');
		 tx_preemp_1t_out	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 tx_preemp_2t	:	IN  STD_LOGIC_VECTOR (4 DOWNTO 0) := (OTHERS => '0');
		 tx_preemp_2t_out	:	OUT  STD_LOGIC_VECTOR (4 DOWNTO 0);
		 tx_vodctrl	:	IN  STD_LOGIC_VECTOR (2 DOWNTO 0) := (OTHERS => '0');
		 tx_vodctrl_out	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0);
		 write_all	:	IN  STD_LOGIC := '0'
	 ); 
 END reconfig_side_alt2gxb_reconfig_4og2;

 ARCHITECTURE RTL OF reconfig_side_alt2gxb_reconfig_4og2 IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF RTL : ARCHITECTURE IS "{-to address_pres_reg[11]} DPRIO_CHANNEL_NUM=11;{-to address_pres_reg[10]} DPRIO_CHANNEL_NUM=10;{-to address_pres_reg[9]} DPRIO_CHANNEL_NUM=9;{-to address_pres_reg[8]} DPRIO_CHANNEL_NUM=8;{-to address_pres_reg[7]} DPRIO_CHANNEL_NUM=7;{-to address_pres_reg[6]} DPRIO_CHANNEL_NUM=6;{-to address_pres_reg[5]} DPRIO_CHANNEL_NUM=5;{-to address_pres_reg[4]} DPRIO_CHANNEL_NUM=4;{-to address_pres_reg[3]} DPRIO_CHANNEL_NUM=3;{-to address_pres_reg[2]} DPRIO_CHANNEL_NUM=2;{-to address_pres_reg[1]} DPRIO_CHANNEL_NUM=1;{-to address_pres_reg[0]} DPRIO_CHANNEL_NUM=0";

	 SIGNAL  wire_calibration_w_lg_w_lg_busy377w428w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy377w391w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy377w378w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_busy392w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_busy379w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_busy377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_busy	:	STD_LOGIC;
	 SIGNAL  wire_calibration_dprio_addr	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_dprio_dataout	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_dprio_rden	:	STD_LOGIC;
	 SIGNAL  wire_calibration_dprio_wren	:	STD_LOGIC;
	 SIGNAL  wire_calibration_quad_addr	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_calibration_reset	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_offset_cancellation_reset207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_calibration_retain_addr	:	STD_LOGIC;
	 SIGNAL  wire_dfe_i_avmm_saddress	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dfe_i_avmm_sread	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_ctrl_read366w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dfe_i_avmm_swrite	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_ctrl_write367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dfe_i_avmm_swritedata	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dfe_i_resetn	:	STD_LOGIC;
	 SIGNAL  wire_dfe_o_avmm_sreaddata	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dfe_o_avmm_swaitrequest	:	STD_LOGIC;
	 SIGNAL  wire_dfe_o_dprio_addr	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dfe_o_dprio_data	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dfe_o_dprio_rden	:	STD_LOGIC;
	 SIGNAL  wire_dfe_o_dprio_wren	:	STD_LOGIC;
	 SIGNAL  wire_dfe_o_quad_address	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_dfe_o_reconfig_busy	:	STD_LOGIC;
	 SIGNAL  wire_dprio_w_lg_w_lg_w_dataout_range1091w1092w1104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range1091w1100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range1091w1095w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range884w1093w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range884w1103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range1075w1076w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_busy567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range1071w1074w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range1094w1099w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range1091w1092w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_w_dataout_range1091w1092w1104w1105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_dataout_range1091w1100w1101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_dataout_range1091w1095w1096w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_lg_w_dataout_range1079w1080w1081w1082w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_lg_w_dataout_range1079w1080w1081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_lg_w_dataout_range1079w1080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_address	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy392w393w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_busy	:	STD_LOGIC;
	 SIGNAL  wire_dprio_datain	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_calibration_w_lg_w_lg_busy379w380w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_dataout	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_dprio_dpriodisable	:	STD_LOGIC;
	 SIGNAL  wire_dprio_dprioin	:	STD_LOGIC;
	 SIGNAL  wire_dprio_dprioload	:	STD_LOGIC;
	 SIGNAL  wire_dprio_rden	:	STD_LOGIC;
	 SIGNAL  wire_calibration_w_lg_w_lg_busy413w414w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_wren	:	STD_LOGIC;
	 SIGNAL  wire_calibration_w_lg_w_lg_busy417w418w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_wren_data	:	STD_LOGIC;
	 SIGNAL  wire_calibration_w_lg_w_lg_busy429w430w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range1071w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range1094w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range1091w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range797w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range884w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range1117w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range1136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range1129w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range1079w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range1075w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range1078w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprio_w_dataout_range1146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_eyemonitor_i_avmm_saddress	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_eyemonitor_i_avmm_sread	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_ctrl_read358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_eyemonitor_i_avmm_swrite	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_ctrl_write359w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_eyemonitor_i_avmm_swritedata	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_eyemonitor_i_resetn	:	STD_LOGIC;
	 SIGNAL  wire_eyemonitor_o_avmm_sreaddata	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_eyemonitor_o_avmm_swaitrequest	:	STD_LOGIC;
	 SIGNAL  wire_eyemonitor_o_dprio_addr	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_eyemonitor_o_dprio_data	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_eyemonitor_o_dprio_rden	:	STD_LOGIC;
	 SIGNAL  wire_eyemonitor_o_dprio_wren	:	STD_LOGIC;
	 SIGNAL  wire_eyemonitor_o_quad_address	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_eyemonitor_o_reconfig_busy	:	STD_LOGIC;
	 SIGNAL	 address_pres_reg	:	STD_LOGIC_VECTOR(11 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF address_pres_reg : SIGNAL IS "PRESERVE_REGISTER=ON";

	 SIGNAL  wire_address_pres_reg_w_lg_w_lg_w_q_range191w192w193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_lg_w_q_range195w196w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_lg_w_q_range191w192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_lg_w_lg_w_lg_w_q_range191w192w193w194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range195w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_w_q_range191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 data_valid_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF data_valid_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_data_valid_reg_ena	:	STD_LOGIC;
	 SIGNAL	 dprio_pulse_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF dprio_pulse_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_dprio_pulse_reg_ena	:	STD_LOGIC;
	 SIGNAL	 error_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 is_illegal_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 reconf_mode_sel_reg	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reconf_mode_sel_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 reset_system_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF reset_system_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_reset_system_reg_sclr	:	STD_LOGIC;
	 SIGNAL	 wire_rx_eqctrl_reg_d	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL	 rx_eqctrl_reg	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rx_eqctrl_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_rx_eqctrl_reg_ena	:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL	 wire_rx_equalizer_dcgain_reg_d	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL	 rx_equalizer_dcgain_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF rx_equalizer_dcgain_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_rx_equalizer_dcgain_reg_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL	 state_mc_reg	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := "00"
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF state_mc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_state_mc_reg_w_lg_q31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_lg_q29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_state_mc_reg_w_q_range67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 tx_preemp_0t_inv_reg	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF tx_preemp_0t_inv_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_tx_preemp_0t_inv_reg_ena	:	STD_LOGIC_VECTOR(0 DOWNTO 0);
	 SIGNAL  wire_tx_preemp_0t_inv_reg_w_lg_w_q_range1139w1140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_preemp_0t_inv_reg_w_q_range1139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 tx_preemp_2t_inv_reg	:	STD_LOGIC_VECTOR(0 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF tx_preemp_2t_inv_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_tx_preemp_2t_inv_reg_ena	:	STD_LOGIC_VECTOR(0 DOWNTO 0);
	 SIGNAL  wire_tx_preemp_2t_inv_reg_w_lg_w_q_range1149w1150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_tx_preemp_2t_inv_reg_w_q_range1149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wire_tx_preemphasisctrl_1stposttap_reg_d	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL	 tx_preemphasisctrl_1stposttap_reg	:	STD_LOGIC_VECTOR(4 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF tx_preemphasisctrl_1stposttap_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_tx_preemphasisctrl_1stposttap_reg_ena	:	STD_LOGIC_VECTOR(4 DOWNTO 0);
	 SIGNAL	 wire_tx_preemphasisctrl_2ndposttap_reg_d	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL	 tx_preemphasisctrl_2ndposttap_reg	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF tx_preemphasisctrl_2ndposttap_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_tx_preemphasisctrl_2ndposttap_reg_ena	:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL	 wire_tx_preemphasisctrl_pretap_reg_d	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL	 tx_preemphasisctrl_pretap_reg	:	STD_LOGIC_VECTOR(3 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF tx_preemphasisctrl_pretap_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_tx_preemphasisctrl_pretap_reg_ena	:	STD_LOGIC_VECTOR(3 DOWNTO 0);
	 SIGNAL	 wire_tx_vodctrl_reg_d	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL	 tx_vodctrl_reg	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF tx_vodctrl_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_tx_vodctrl_reg_ena	:	STD_LOGIC_VECTOR(2 DOWNTO 0);
	 SIGNAL	 wr_addr_inc_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_addr_inc_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wr_rd_pulse_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wr_rd_pulse_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_wr_rd_pulse_reg_ena	:	STD_LOGIC;
	 SIGNAL	 wire_wr_rd_pulse_reg_sclr	:	STD_LOGIC;
	 SIGNAL  wire_wr_rd_pulse_reg_w_lg_q617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wr_rd_pulse_reg_w_lg_q570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 wren_data_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF wren_data_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL	 wire_wren_data_reg_ena	:	STD_LOGIC;
	 SIGNAL  wire_wren_data_reg_w_lg_w_lg_q724w725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wren_data_reg_w_lg_q723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wren_data_reg_w_lg_q724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_wren_data_reg_w_lg_q728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub1_dataa	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub11_add_sub	:	STD_LOGIC;
	 SIGNAL  wire_add_sub11_dataa	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub11_result	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub12_add_sub	:	STD_LOGIC;
	 SIGNAL  wire_add_sub12_dataa	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub12_result	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub2_dataa	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub2_result	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cmpr10_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr10_datab	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cmpr7_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr7_datab	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cmpr8_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr8_datab	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_cmpr9_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr9_datab	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_max_oper_limit_w_lg_aeb118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_max_oper_limit_aeb	:	STD_LOGIC;
	 SIGNAL  wire_gnd	:	STD_LOGIC;
	 SIGNAL  wire_addr_cntr_q	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_addr_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_write_done623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_addr_cntr_sload	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_idle_state625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_oper_count_q	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_oper_count_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_idle_state102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_w_lg_w_q_range695w698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_w_lg_w_q_range693w696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_w_lg_w_q_range693w708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_w_lg_w_q_range699w700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_cnt_en	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_read_addr_inc674w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_data	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_read_done675w676w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_sload	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_idle_state683w684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_w_q_range695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_w_q_range699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_read_addr_cntr_w_q_range693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_lg_w_q_range930w933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_lg_w_q_range928w951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_lg_w_q_range928w931w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_lg_w_q_range934w943w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_lg_w_q_range934w935w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_data	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_q	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_sclr	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_write_done910w911w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_sload	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_idle_state918w919w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_q_range930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_q_range934w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_write_addr_cntr_w_q_range928w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_chl_addr_decode_eq	:	STD_LOGIC_VECTOR (143 DOWNTO 0);
	 SIGNAL  wire_reconf_mode_dec_eq	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_adce_dprio_addr_mux_data	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_adce_dprio_addr_mux_result	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_adce_dprio_addr_mux_sel	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_adce_dprio_data_mux_data	:	STD_LOGIC_VECTOR (63 DOWNTO 0);
	 SIGNAL  wire_adce_dprio_data_mux_result	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_adce_dprio_data_mux_sel	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_adce_dprio_enas_mux_data	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_adce_dprio_enas_mux_result	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_adce_dprio_enas_mux_sel	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_mux_data	:	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_mux_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_address_pres_reg_mux_sel	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_aeq_ch_done_mux_result	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprioout_mux_result	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_dprioout_mux_sel	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_s2_to_058w59w60w61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_s2_to_058w70w71w72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range842w843w844w867w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range842w846w860w861w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w876w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_header_proc593w594w595w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_s2_to_058w59w60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_s2_to_058w70w71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range842w850w851w852w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w1021w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dprio_datain735w736w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_analog_control108w109w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_analog_control106w107w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1613w615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_gt_0_964w996w1000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_word_done906w907w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range840w848w849w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range840w871w872w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range842w843w844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range842w869w870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range842w846w868w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range842w846w860w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range842w846w847w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1033w1034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1022w1023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range842w873w874w875w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_adce_busy_state132w133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_adce_busy_state132w448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_adce_busy_state132w461w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_adce_busy_state132w473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_adce_busy_state132w485w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_adce_busy_state132w497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_adce_busy_state132w509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy182w183w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy182w511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy182w520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy182w528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy182w536w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy182w544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy182w552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_header_proc593w594w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_bonded_global_clk_div9w10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_bonded_reconfig17w18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_table_3313w14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_s2_to_058w59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_s2_to_058w70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_tx_reconfig93w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range842w850w851w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv959w_range1011w1018w1043w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv959w_range1011w1018w1054w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1019w1020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w156w157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w752w753w754w755w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_tier_1737w738w739w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dprio_datain_68_6B742w743w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mif_type_error95w96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_channel_address_range153w154w155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_channel_address_range143w144w145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_logical_pll_sel_num_range150w151w152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_logical_pll_sel_num_range139w140w141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_adce_busy_state444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_adce_busy_state458w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_adce_busy_state470w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_adce_busy_state482w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_adce_busy_state494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_adce_busy_state506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy186w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_ctrl_address357w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_ctrl_address365w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_ctrl_writedata360w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_ctrl_writedata368w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dfe_busy436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dfe_busy452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dfe_busy464w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dfe_busy476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dfe_busy488w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dfe_busy500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain735w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_64_67744w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_7c_7f741w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_7c_7f_inv740w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_preemp1t747w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_vodctrl749w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_pulse709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_pulse716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_eyemon_busy440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_eyemon_busy455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_eyemon_busy467w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_eyemon_busy479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_eyemon_busy491w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_eyemon_busy503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_adce_mode_sel103w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_analog_control108w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_analog_control106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_bonded_reconfig23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_bonded_reconfig16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_illegal_reg_d124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_illegal_reg_out121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_3312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_59138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_61148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1589w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1105w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tx_local_div_ctrl104w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_w_lg_read49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_address560w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state1114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state1068w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state1088w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state1111w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state1124w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state1118w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state1147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state1137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state1130w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_word_64_67_data_valid1085w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_word_68_6B_data_valid1065w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_word_7c_7f_data_valid1126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_word_7c_7f_inv_data_valid703w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_word_preemp_1t_data_valid1121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_word_vodctrl_data_valid1108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_eq_0_1004w1060w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_eq_10_1045w1057w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_eq_3_1026w1059w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_eq_6_1036w1058w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_gt_0_964w992w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_gt_0_964w996w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_wr_pulse732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_wr_pulse729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_address561w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_all25w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state1135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state1145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state1067w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state1087w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state1123w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state1110w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state1084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state1064w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state1113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state1120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state1107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state1116w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state1128w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_word_7c_7f_inv_data_valid938w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_word_done906w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_reconfig_mode_sel_range644w645w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range838w854w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range838w864w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range840w848w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range840w871w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range842w843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range842w869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range842w846w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqdcgain_range820w821w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_vodctrl_range761w769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_vodctrl_range761w762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_vodctrl_range759w771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_vodctrl_range759w763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv959w_range1014w1015w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv959w_range1014w1033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv959w_range1014w1022w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_done120w123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range842w873w874w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_tx_vodctrl_range759w760w768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv959w_range1011w1012w1013w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1041w1042w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_adce_busy_state132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bonded_skip604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_cal_busy182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_pulse581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_header_proc593w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_idle_state117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_adce116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_analog_control731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_bonded_global_clk_div9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_bonded_reconfig17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_central_pcs149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_cruclk_addr0606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_diff_mif564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_do_dfe356w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_do_eyemon364w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_global_clk_div_mode602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_illegal_reg_d579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_illegal_reg_out122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_pll_address142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_protected_bit603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rcxpat_chnl_en_ch607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_table_3313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rd_pulse198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_done580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_state571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reconfig_reset_all28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reset_reconf_addr592w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rx_reconfig92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s0_to_056w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s0_to_157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s1_to_068w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s1_to_169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s2_to_058w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_tx_reconfig93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_gt_10_982w989w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_gt_3_970w991w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_gt_6_976w990w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_wr_pulse199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_all_int47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_done91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_skip605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_state48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_reconfig_mode_sel_range85w643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range845w853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range838w839w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range840w841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range842w850w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_preemp_0t_range2w896w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_preemp_2t_range4w900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_vodctrl_range758w770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv959w_range1010w1017w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv959w_range1011w1018w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv959w_range1014w1019w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w876w877w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w1024w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_cal_busy182w511w512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_cal_busy182w520w521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_cal_busy182w528w529w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_cal_busy182w536w537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_cal_busy182w544w545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_cal_busy182w552w553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_bonded_global_clk_div9w10w11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_table_3313w14w15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w1052w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w1055w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w156w157w158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_mif_type_error95w96w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy186w187w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy516w517w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy525w526w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy533w534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy541w542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy549w550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_cal_busy557w558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dprio_datain_vodctrl749w750w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_state1114w1115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_state1068w1069w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_state1088w1089w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_state1111w1112w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_state1124w1125w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_state1118w1119w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_state1130w1131w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_word_64_67_data_valid1085w1086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_word_68_6B_data_valid1065w1066w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_word_7c_7f_data_valid1126w1127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_word_preemp_1t_data_valid1121w1122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_read_word_vodctrl_data_valid1108w1109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range838w854w855w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqctrl_range838w864w865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_tx_vodctrl_range759w771w772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_tx_vodctrl_range759w763w764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_bonded_reconfig17w24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1590w616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1590w591w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w876w877w878w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w511w512w513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w520w521w522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w528w529w530w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w536w537w538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w544w545w546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w552w553w554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_mif_type_error95w96w97w98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w146w147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_dprio_datain_vodctrl749w750w751w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range838w854w855w856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w876w877w878w879w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w514w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w752w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w857w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_w_lg_w876w877w878w879w880w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w752w753w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w857w858w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w752w753w754w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_w587w588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch584w585w586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_adce39w40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_pll_address135w136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_rcxpat_chnl_en_ch584w585w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_is_tier_1737w738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_s0_to_262w63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_s0_to_273w74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_write_word_preemp1t_data_valid745w746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_rx_eqdcgain_range816w824w826w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1049w1050w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_adce_busy_state128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dprio_datain_68_6B742w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_adce39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_do_eyemon131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_pll_address135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_rcxpat_chnl_en_ch584w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_is_tier_1737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mif_type_error95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_read_done120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_reset_system575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s0_to_262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_s0_to_273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_word_preemp1t_data_valid745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_write_word_vodctrl_data_valid748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_channel_address_range153w154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_channel_address_range143w144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_logical_pll_sel_num_range150w151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_logical_pll_sel_num_range139w140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqdcgain_range816w822w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqdcgain_range816w824w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv959w_range1014w1049w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range845w863w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range840w862w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_rx_eqctrl_range842w873w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_tx_vodctrl_range759w760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv959w_range1011w1012w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_w_rx_eqv959w_range1014w1041w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  a2gr_dprio_addr :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  a2gr_dprio_data :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  a2gr_dprio_rden :	STD_LOGIC;
	 SIGNAL  a2gr_dprio_wren :	STD_LOGIC;
	 SIGNAL  a2gr_dprio_wren_data :	STD_LOGIC;
	 SIGNAL  adce_busy_state :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  adce_dprio_addr_s4 :	STD_LOGIC_VECTOR (15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  adce_dprio_data :	STD_LOGIC_VECTOR (15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  adce_dprio_rden :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  adce_dprio_wren :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  adce_error_wire :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  adce_pres_reg :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  adce_quad_addr_s4 :	STD_LOGIC_VECTOR (8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  adce_state :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  aeq_ch_done :	STD_LOGIC_VECTOR (143 DOWNTO 0);
	 SIGNAL  analog_read_max_limit :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  analog_write_max_limit :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  bonded_skip :	STD_LOGIC;
	 SIGNAL  busy_state :	STD_LOGIC;
	 SIGNAL  cal_busy :	STD_LOGIC;
	 SIGNAL  cal_channel_address :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  cal_channel_address_out :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  cal_dprio_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  cal_dprioout_wire :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  cal_quad_address :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  cal_testbuses :	STD_LOGIC_VECTOR (575 DOWNTO 0);
	 SIGNAL  channel_address :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  channel_address_out :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  default_max_limit_wire :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  dfe_busy :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  dfe_dprio_addr :	STD_LOGIC_VECTOR (15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  dfe_dprio_data :	STD_LOGIC_VECTOR (15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  dfe_dprio_rden :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  dfe_dprio_wren :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  dfe_pres_reg :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  dfe_quad_address :	STD_LOGIC_VECTOR (8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  dfe_readdata :	STD_LOGIC_VECTOR (15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  dfe_swaitrequest :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  diff_mif_wr_rd_busy :	STD_LOGIC;
	 SIGNAL  dprio_datain :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_64_67 :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_68_6B :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_7c_7f :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_7c_7f_inv :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_preemp1t :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_datain_vodctrl :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  dprio_pulse :	STD_LOGIC;
	 SIGNAL  en_read_trigger :	STD_LOGIC
	 -- synopsys translate_off
	  := '1'
	 -- synopsys translate_on
	 ;
	 SIGNAL  en_write_trigger :	STD_LOGIC
	 -- synopsys translate_off
	  := '1'
	 -- synopsys translate_on
	 ;
	 SIGNAL  eyemon_busy :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  eyemon_dprio_addr :	STD_LOGIC_VECTOR (15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  eyemon_dprio_data :	STD_LOGIC_VECTOR (15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  eyemon_dprio_rden :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  eyemon_dprio_wren :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  eyemon_pres_reg :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  eyemon_quad_address :	STD_LOGIC_VECTOR (8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  eyemon_readdata :	STD_LOGIC_VECTOR (15 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  eyemon_swaitrequest :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  header_proc :	STD_LOGIC;
	 SIGNAL  idle_state :	STD_LOGIC;
	 SIGNAL  internal_write_pulse :	STD_LOGIC;
	 SIGNAL  invalid_eq_dcgain :	STD_LOGIC;
	 SIGNAL  is_adce :	STD_LOGIC;
	 SIGNAL  is_adce_all_control :	STD_LOGIC;
	 SIGNAL  is_adce_continuous_single_control :	STD_LOGIC;
	 SIGNAL  is_adce_mode_sel :	STD_LOGIC;
	 SIGNAL  is_adce_one_time_single_control :	STD_LOGIC;
	 SIGNAL  is_adce_single_control :	STD_LOGIC;
	 SIGNAL  is_adce_standby_single_control :	STD_LOGIC;
	 SIGNAL  is_analog_control :	STD_LOGIC;
	 SIGNAL  is_bonded_global_clk_div :	STD_LOGIC;
	 SIGNAL  is_bonded_reconfig :	STD_LOGIC;
	 SIGNAL  is_central_pcs :	STD_LOGIC;
	 SIGNAL  is_cruclk_addr0 :	STD_LOGIC;
	 SIGNAL  is_diff_mif :	STD_LOGIC;
	 SIGNAL  is_do_dfe :	STD_LOGIC;
	 SIGNAL  is_do_eyemon :	STD_LOGIC;
	 SIGNAL  is_global_clk_div_mode :	STD_LOGIC;
	 SIGNAL  is_illegal_reg_d :	STD_LOGIC;
	 SIGNAL  is_illegal_reg_out :	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  is_pll_address :	STD_LOGIC;
	 SIGNAL  is_protected_bit :	STD_LOGIC;
	 SIGNAL  is_rcxpat_chnl_en_ch :	STD_LOGIC;
	 SIGNAL  is_table_33 :	STD_LOGIC;
	 SIGNAL  is_table_59 :	STD_LOGIC;
	 SIGNAL  is_table_61 :	STD_LOGIC;
	 SIGNAL  is_tier_1 :	STD_LOGIC;
	 SIGNAL  is_tier_2 :	STD_LOGIC;
	 SIGNAL  is_tx_local_div_ctrl :	STD_LOGIC;
	 SIGNAL  local_ch_dec :	STD_LOGIC;
	 SIGNAL  logical_pll_sel_num :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  mif_family_error :	STD_LOGIC;
	 SIGNAL  mif_reconfig_done :	STD_LOGIC;
	 SIGNAL  mif_type_error :	STD_LOGIC;
	 SIGNAL  offset_cancellation_reset	:	STD_LOGIC;
	 SIGNAL  quad_address :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  quad_address_out :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  rate_switch_ctrl_max_limit :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  rd_pulse :	STD_LOGIC;
	 SIGNAL  read_addr_inc :	STD_LOGIC;
	 SIGNAL  read_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  read_done :	STD_LOGIC;
	 SIGNAL  read_state :	STD_LOGIC;
	 SIGNAL  read_word_64_67_data_valid :	STD_LOGIC;
	 SIGNAL  read_word_68_6B_data_valid :	STD_LOGIC;
	 SIGNAL  read_word_7c_7f_data_valid :	STD_LOGIC;
	 SIGNAL  read_word_7c_7f_inv_data_valid :	STD_LOGIC;
	 SIGNAL  read_word_done :	STD_LOGIC;
	 SIGNAL  read_word_preemp_1t_data_valid :	STD_LOGIC;
	 SIGNAL  read_word_vodctrl_data_valid :	STD_LOGIC;
	 SIGNAL  reconfig_datain :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  reconfig_reset_all :	STD_LOGIC;
	 SIGNAL  remap_eyemon :	STD_LOGIC;
	 SIGNAL  reset_addr_done :	STD_LOGIC;
	 SIGNAL  reset_reconf_addr :	STD_LOGIC;
	 SIGNAL  reset_system :	STD_LOGIC;
	 SIGNAL  rx_reconfig :	STD_LOGIC;
	 SIGNAL  s0_to_0 :	STD_LOGIC;
	 SIGNAL  s0_to_1 :	STD_LOGIC;
	 SIGNAL  s0_to_2 :	STD_LOGIC;
	 SIGNAL  s1_to_0 :	STD_LOGIC;
	 SIGNAL  s1_to_1 :	STD_LOGIC;
	 SIGNAL  s2_to_0 :	STD_LOGIC;
	 SIGNAL  sel_max_limit :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  start	:	STD_LOGIC;
	 SIGNAL  state_mc_reg_in :	STD_LOGIC_VECTOR (1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  tier_1_max_limit :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  transceiver_init	:	STD_LOGIC;
	 SIGNAL  tx_preemp_0t_out_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_preemp_0t_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_preemp_2t_out_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_preemp_2t_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  tx_reconfig :	STD_LOGIC;
	 SIGNAL  wire_w185w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  w721w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  w_eq_0_1004w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_eq_10_1045w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_eq_3_1026w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_eq_6_1036w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_gt_0_964w :	STD_LOGIC;
	 SIGNAL  w_gt_0_only988w :	STD_LOGIC;
	 SIGNAL  w_gt_10_982w :	STD_LOGIC;
	 SIGNAL  w_gt_10_only1002w :	STD_LOGIC;
	 SIGNAL  w_gt_3_970w :	STD_LOGIC;
	 SIGNAL  w_gt_3_only995w :	STD_LOGIC;
	 SIGNAL  w_gt_6_976w :	STD_LOGIC;
	 SIGNAL  w_gt_6_only999w :	STD_LOGIC;
	 SIGNAL  w_rx_eqa958w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  w_rx_eqb957w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  w_rx_eqc956w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  w_rx_eqctrl_out954w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  w_rx_eqd955w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  w_rx_eqdcgain_out1070w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  w_rx_eqv959w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  w_tx_vodctrl_out1090w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  w_wire_adce_dprioout_mux2434w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  w_wire_adce_dprioout_mux433w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  w_wire_dfe_dprioout_mux431w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  w_wire_eyemon_dprioout_mux432w :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wr_pulse :	STD_LOGIC;
	 SIGNAL  write_addr_inc :	STD_LOGIC;
	 SIGNAL  write_address :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  write_all_int :	STD_LOGIC;
	 SIGNAL  write_done :	STD_LOGIC;
	 SIGNAL  write_happened :	STD_LOGIC;
	 SIGNAL  write_skip :	STD_LOGIC;
	 SIGNAL  write_state :	STD_LOGIC;
	 SIGNAL  write_word_64_67_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_68_6B_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_7c_7f_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_7c_7f_inv_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_done :	STD_LOGIC;
	 SIGNAL  write_word_preemp1t_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_preemp1ta_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_preemp1tb_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_vodctrl_data_valid :	STD_LOGIC;
	 SIGNAL  write_word_vodctrla_data_valid :	STD_LOGIC;
	 SIGNAL  wire_w_adce_quad_addr_s4_range443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_adce_quad_addr_s4_range457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_adce_quad_addr_s4_range469w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_adce_quad_addr_s4_range481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_adce_quad_addr_s4_range493w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_adce_quad_addr_s4_range505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_cal_quad_address_range515w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_cal_quad_address_range524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_cal_quad_address_range532w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_cal_quad_address_range540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_cal_quad_address_range548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_cal_quad_address_range556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_range153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_channel_address_range143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dfe_quad_address_range435w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dfe_quad_address_range451w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dfe_quad_address_range463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dfe_quad_address_range475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dfe_quad_address_range487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_dfe_quad_address_range499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_eyemon_quad_address_range439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_eyemon_quad_address_range454w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_eyemon_quad_address_range466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_eyemon_quad_address_range478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_eyemon_quad_address_range490w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_eyemon_quad_address_range502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_logical_pll_sel_num_range150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_logical_pll_sel_num_range139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_quad_address_range447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_quad_address_range460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_quad_address_range472w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_quad_address_range484w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_quad_address_range496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_quad_address_range508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_reconfig_mode_sel_range644w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_reconfig_mode_sel_range85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_eqctrl_range845w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_eqctrl_range838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_eqctrl_range840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_eqctrl_range842w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_eqdcgain_range819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_eqdcgain_range820w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_rx_eqdcgain_range816w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tx_preemp_0t_range2w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tx_preemp_0t_wire_range894w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_tx_preemp_2t_range4w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tx_preemp_2t_wire_range898w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_w_tx_vodctrl_range761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tx_vodctrl_range758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_tx_vodctrl_range759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_rx_eqv959w_range1010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_rx_eqv959w_range1011w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_rx_eqv959w_range1014w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_adce_dprioout_mux2434w_range449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_adce_dprioout_mux2434w_range462w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_adce_dprioout_mux2434w_range474w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_adce_dprioout_mux2434w_range486w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_adce_dprioout_mux2434w_range498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_adce_dprioout_mux2434w_range510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_adce_dprioout_mux433w_range445w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_adce_dprioout_mux433w_range459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_adce_dprioout_mux433w_range471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_adce_dprioout_mux433w_range483w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_adce_dprioout_mux433w_range495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_adce_dprioout_mux433w_range507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_dfe_dprioout_mux431w_range437w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_dfe_dprioout_mux431w_range453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_dfe_dprioout_mux431w_range465w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_dfe_dprioout_mux431w_range477w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_dfe_dprioout_mux431w_range489w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_dfe_dprioout_mux431w_range501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_eyemon_dprioout_mux432w_range441w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_eyemon_dprioout_mux432w_range456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_eyemon_dprioout_mux432w_range468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_eyemon_dprioout_mux432w_range480w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_eyemon_dprioout_mux432w_range492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_w_wire_eyemon_dprioout_mux432w_range504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  alt_cal
	 GENERIC 
	 (
		CHANNEL_ADDRESS_WIDTH	:	NATURAL := 1;
		NUMBER_OF_CHANNELS	:	NATURAL;
		SIM_MODEL_MODE	:	STRING := "FALSE";
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "alt_cal"
	 );
	 PORT
	 ( 
		busy	:	OUT STD_LOGIC;
		cal_error	:	OUT STD_LOGIC_VECTOR(NUMBER_OF_CHANNELS-1 DOWNTO 0);
		clock	:	IN STD_LOGIC;
		dprio_addr	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_busy	:	IN STD_LOGIC;
		dprio_datain	:	IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_dataout	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		dprio_rden	:	OUT STD_LOGIC;
		dprio_wren	:	OUT STD_LOGIC;
		quad_addr	:	OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		remap_addr	:	IN STD_LOGIC_VECTOR(11 DOWNTO 0) := (OTHERS => '0');
		reset	:	IN STD_LOGIC := '0';
		retain_addr	:	OUT STD_LOGIC;
		start	:	IN STD_LOGIC := '0';
		testbuses	:	IN STD_LOGIC_VECTOR(NUMBER_OF_CHANNELS*4-1 DOWNTO 0) := (OTHERS => '0');
		transceiver_init	:	IN STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  alt_dfe
	 GENERIC 
	 (
		avmm_master_addr_width	:	NATURAL := 16;
		avmm_master_rdata_width	:	NATURAL := 16;
		avmm_master_wdata_width	:	NATURAL := 16;
		avmm_slave_addr_width	:	NATURAL := 16;
		avmm_slave_rdata_width	:	NATURAL := 16;
		avmm_slave_wdata_width	:	NATURAL := 16;
		channel_address_width	:	NATURAL;
		dprio_addr_width	:	NATURAL := 16;
		dprio_data_width	:	NATURAL := 16;
		ireg_chaddr_width	:	NATURAL;
		ireg_data_width	:	NATURAL := 16;
		ireg_wdaddr_width	:	NATURAL := 2;
		lpm_type	:	STRING := "alt_dfe"
	 );
	 PORT
	 ( 
		i_avmm_clk	:	IN STD_LOGIC;
		i_avmm_saddress	:	IN STD_LOGIC_VECTOR(avmm_slave_addr_width-1 DOWNTO 0);
		i_avmm_sread	:	IN STD_LOGIC;
		i_avmm_swrite	:	IN STD_LOGIC;
		i_avmm_swritedata	:	IN STD_LOGIC_VECTOR(avmm_slave_wdata_width-1 DOWNTO 0);
		i_dprio_busy	:	IN STD_LOGIC;
		i_dprio_in	:	IN STD_LOGIC_VECTOR(dprio_data_width-1 DOWNTO 0);
		i_remap_address	:	IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		i_resetn	:	IN STD_LOGIC;
		o_avmm_sreaddata	:	OUT STD_LOGIC_VECTOR(avmm_slave_rdata_width-1 DOWNTO 0);
		o_avmm_swaitrequest	:	OUT STD_LOGIC;
		o_dprio_addr	:	OUT STD_LOGIC_VECTOR(dprio_addr_width-1 DOWNTO 0);
		o_dprio_data	:	OUT STD_LOGIC_VECTOR(dprio_data_width-1 DOWNTO 0);
		o_dprio_rden	:	OUT STD_LOGIC;
		o_dprio_wren	:	OUT STD_LOGIC;
		o_quad_address	:	OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		o_reconfig_busy	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  reconfig_side_alt_dprio_2vj
	 PORT
	 ( 
		address	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0);
		busy	:	OUT  STD_LOGIC;
		datain	:	IN  STD_LOGIC_VECTOR(15 DOWNTO 0) := (OTHERS => '0');
		dataout	:	OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		dpclk	:	IN  STD_LOGIC;
		dpriodisable	:	OUT  STD_LOGIC;
		dprioin	:	OUT  STD_LOGIC;
		dprioload	:	OUT  STD_LOGIC;
		dprioout	:	IN  STD_LOGIC;
		quad_address	:	IN  STD_LOGIC_VECTOR(8 DOWNTO 0);
		rden	:	IN  STD_LOGIC := '0';
		reset	:	IN  STD_LOGIC := '0';
		wren	:	IN  STD_LOGIC := '0';
		wren_data	:	IN  STD_LOGIC := '0'
	 ); 
	 END COMPONENT;
	 COMPONENT  alt_eyemon
	 GENERIC 
	 (
		avmm_master_addr_width	:	NATURAL := 16;
		avmm_master_rdata_width	:	NATURAL := 16;
		avmm_master_wdata_width	:	NATURAL := 16;
		avmm_slave_addr_width	:	NATURAL := 16;
		avmm_slave_rdata_width	:	NATURAL := 16;
		avmm_slave_wdata_width	:	NATURAL := 16;
		channel_address_width	:	NATURAL;
		dprio_addr_width	:	NATURAL := 16;
		dprio_data_width	:	NATURAL := 16;
		ireg_chaddr_width	:	NATURAL;
		ireg_data_width	:	NATURAL := 16;
		ireg_wdaddr_width	:	NATURAL := 2;
		lpm_type	:	STRING := "alt_eyemon"
	 );
	 PORT
	 ( 
		i_avmm_clk	:	IN STD_LOGIC;
		i_avmm_saddress	:	IN STD_LOGIC_VECTOR(avmm_slave_addr_width-1 DOWNTO 0);
		i_avmm_sread	:	IN STD_LOGIC;
		i_avmm_swrite	:	IN STD_LOGIC;
		i_avmm_swritedata	:	IN STD_LOGIC_VECTOR(avmm_slave_wdata_width-1 DOWNTO 0);
		i_dprio_busy	:	IN STD_LOGIC;
		i_dprio_in	:	IN STD_LOGIC_VECTOR(dprio_data_width-1 DOWNTO 0);
		i_remap_address	:	IN STD_LOGIC_VECTOR(11 DOWNTO 0);
		i_remap_phase	:	IN STD_LOGIC;
		i_resetn	:	IN STD_LOGIC;
		o_avmm_sreaddata	:	OUT STD_LOGIC_VECTOR(avmm_slave_rdata_width-1 DOWNTO 0);
		o_avmm_swaitrequest	:	OUT STD_LOGIC;
		o_dprio_addr	:	OUT STD_LOGIC_VECTOR(dprio_addr_width-1 DOWNTO 0);
		o_dprio_data	:	OUT STD_LOGIC_VECTOR(dprio_data_width-1 DOWNTO 0);
		o_dprio_rden	:	OUT STD_LOGIC;
		o_dprio_wren	:	OUT STD_LOGIC;
		o_quad_address	:	OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
		o_reconfig_busy	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_counter
	 GENERIC 
	 (
		lpm_avalue	:	STRING := "0";
		lpm_direction	:	STRING := "DEFAULT";
		lpm_modulus	:	NATURAL := 0;
		lpm_port_updown	:	STRING := "PORT_CONNECTIVITY";
		lpm_pvalue	:	STRING := "0";
		lpm_svalue	:	STRING := "0";
		lpm_width	:	NATURAL;
		lpm_type	:	STRING := "lpm_counter"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aload	:	IN STD_LOGIC := '0';
		aset	:	IN STD_LOGIC := '0';
		cin	:	IN STD_LOGIC := '1';
		clk_en	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC;
		cnt_en	:	IN STD_LOGIC := '1';
		cout	:	OUT STD_LOGIC;
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		eq	:	OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		q	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0);
		sclr	:	IN STD_LOGIC := '0';
		sload	:	IN STD_LOGIC := '0';
		sset	:	IN STD_LOGIC := '0';
		updown	:	IN STD_LOGIC := '1'
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_decode
	 GENERIC 
	 (
		LPM_DECODES	:	NATURAL;
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_decode"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		data	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		enable	:	IN STD_LOGIC := '1';
		eq	:	OUT STD_LOGIC_VECTOR(LPM_DECODES-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  reconfig_side_mux_t7a
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(63 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(15 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  reconfig_side_mux_86a
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(1 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  reconfig_side_mux_p7a
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(47 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(11 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  reconfig_side_mux_i9a
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(143 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
	 COMPONENT  reconfig_side_mux_08a
	 PORT
	 ( 
		data	:	IN  STD_LOGIC_VECTOR(35 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(0 DOWNTO 0);
		sel	:	IN  STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_gnd <= '0';
	wire_w_lg_w_lg_w_lg_w_lg_s2_to_058w59w60w61w(0) <= wire_w_lg_w_lg_w_lg_s2_to_058w59w60w(0) AND wire_state_mc_reg_w_q_range55w(0);
	wire_w_lg_w_lg_w_lg_w_lg_s2_to_058w70w71w72w(0) <= wire_w_lg_w_lg_w_lg_s2_to_058w70w71w(0) AND wire_state_mc_reg_w_q_range67w(0);
	wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range842w843w844w867w(0) <= wire_w_lg_w_lg_w_rx_eqctrl_range842w843w844w(0) AND wire_w_rx_eqctrl_range845w(0);
	wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range842w846w860w861w(0) <= wire_w_lg_w_lg_w_rx_eqctrl_range842w846w860w(0) AND wire_w_lg_w_rx_eqctrl_range845w853w(0);
	wire_w876w(0) <= wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range842w873w874w875w(0) AND wire_w_rx_eqctrl_range845w(0);
	wire_w_lg_w_lg_w_lg_header_proc593w594w595w(0) <= wire_w_lg_w_lg_header_proc593w594w(0) AND wire_w_lg_w_lg_is_tier_1590w591w(0);
	wire_w_lg_w_lg_w_lg_s2_to_058w59w60w(0) <= wire_w_lg_w_lg_s2_to_058w59w(0) AND wire_w_lg_s0_to_056w(0);
	wire_w_lg_w_lg_w_lg_s2_to_058w70w71w(0) <= wire_w_lg_w_lg_s2_to_058w70w(0) AND wire_w_lg_s1_to_068w(0);
	wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range842w850w851w852w(0) <= wire_w_lg_w_lg_w_rx_eqctrl_range842w850w851w(0) AND wire_w_rx_eqctrl_range838w(0);
	wire_w1021w(0) <= wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1019w1020w(0) AND wire_w_lg_w_w_rx_eqv959w_range1010w1017w(0);
	loop1 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_dprio_datain735w736w(i) <= wire_w_lg_dprio_datain735w(i) AND write_state;
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 11 GENERATE 
		wire_w_lg_w_lg_is_analog_control108w109w(i) <= wire_w_lg_is_analog_control108w(i) AND write_state;
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 11 GENERATE 
		wire_w_lg_w_lg_is_analog_control106w107w(i) <= wire_w_lg_is_analog_control106w(0) AND analog_read_max_limit(i);
	END GENERATE loop3;
	wire_w_lg_w_lg_is_tier_1613w615w(0) <= wire_w_lg_is_tier_1613w(0) AND wire_w_lg_w587w588w(0);
	wire_w_lg_w_lg_w_gt_0_964w996w1000w(0) <= wire_w_lg_w_gt_0_964w996w(0) AND w_gt_6_976w;
	wire_w_lg_w_lg_write_word_done906w907w(0) <= wire_w_lg_write_word_done906w(0) AND write_happened;
	wire_w_lg_w_lg_w_rx_eqctrl_range840w848w849w(0) <= wire_w_lg_w_rx_eqctrl_range840w848w(0) AND wire_w_rx_eqctrl_range845w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range840w871w872w(0) <= wire_w_lg_w_rx_eqctrl_range840w871w(0) AND wire_w_lg_w_rx_eqctrl_range845w853w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range842w843w844w(0) <= wire_w_lg_w_rx_eqctrl_range842w843w(0) AND wire_w_lg_w_rx_eqctrl_range838w839w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range842w869w870w(0) <= wire_w_lg_w_rx_eqctrl_range842w869w(0) AND wire_w_lg_w_rx_eqctrl_range845w853w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range842w846w868w(0) <= wire_w_lg_w_rx_eqctrl_range842w846w(0) AND wire_w_lg_w_rx_eqctrl_range845w853w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range842w846w860w(0) <= wire_w_lg_w_rx_eqctrl_range842w846w(0) AND wire_w_lg_w_rx_eqctrl_range838w839w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range842w846w847w(0) <= wire_w_lg_w_rx_eqctrl_range842w846w(0) AND wire_w_rx_eqctrl_range845w(0);
	wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1033w1034w(0) <= wire_w_lg_w_w_rx_eqv959w_range1014w1033w(0) AND wire_w_lg_w_w_rx_eqv959w_range1010w1017w(0);
	wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1022w1023w(0) <= wire_w_lg_w_w_rx_eqv959w_range1014w1022w(0) AND wire_w_w_rx_eqv959w_range1010w(0);
	wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range842w873w874w875w(0) <= wire_w_lg_w_lg_w_rx_eqctrl_range842w873w874w(0) AND wire_w_rx_eqctrl_range838w(0);
	wire_w_lg_w_lg_adce_busy_state132w133w(0) <= wire_w_lg_adce_busy_state132w(0) AND wire_w_lg_is_do_eyemon131w(0);
	wire_w_lg_w_lg_adce_busy_state132w448w(0) <= wire_w_lg_adce_busy_state132w(0) AND wire_w_quad_address_range447w(0);
	wire_w_lg_w_lg_adce_busy_state132w461w(0) <= wire_w_lg_adce_busy_state132w(0) AND wire_w_quad_address_range460w(0);
	wire_w_lg_w_lg_adce_busy_state132w473w(0) <= wire_w_lg_adce_busy_state132w(0) AND wire_w_quad_address_range472w(0);
	wire_w_lg_w_lg_adce_busy_state132w485w(0) <= wire_w_lg_adce_busy_state132w(0) AND wire_w_quad_address_range484w(0);
	wire_w_lg_w_lg_adce_busy_state132w497w(0) <= wire_w_lg_adce_busy_state132w(0) AND wire_w_quad_address_range496w(0);
	wire_w_lg_w_lg_adce_busy_state132w509w(0) <= wire_w_lg_adce_busy_state132w(0) AND wire_w_quad_address_range508w(0);
	loop4 : FOR i IN 0 TO 11 GENERATE 
		wire_w_lg_w_lg_cal_busy182w183w(i) <= wire_w_lg_cal_busy182w(0) AND wire_address_pres_reg_mux_result(i);
	END GENERATE loop4;
	wire_w_lg_w_lg_cal_busy182w511w(0) <= wire_w_lg_cal_busy182w(0) AND wire_w_w_wire_dfe_dprioout_mux431w_range437w(0);
	wire_w_lg_w_lg_cal_busy182w520w(0) <= wire_w_lg_cal_busy182w(0) AND wire_w_w_wire_dfe_dprioout_mux431w_range453w(0);
	wire_w_lg_w_lg_cal_busy182w528w(0) <= wire_w_lg_cal_busy182w(0) AND wire_w_w_wire_dfe_dprioout_mux431w_range465w(0);
	wire_w_lg_w_lg_cal_busy182w536w(0) <= wire_w_lg_cal_busy182w(0) AND wire_w_w_wire_dfe_dprioout_mux431w_range477w(0);
	wire_w_lg_w_lg_cal_busy182w544w(0) <= wire_w_lg_cal_busy182w(0) AND wire_w_w_wire_dfe_dprioout_mux431w_range489w(0);
	wire_w_lg_w_lg_cal_busy182w552w(0) <= wire_w_lg_cal_busy182w(0) AND wire_w_w_wire_dfe_dprioout_mux431w_range501w(0);
	wire_w_lg_w_lg_header_proc593w594w(0) <= wire_w_lg_header_proc593w(0) AND wire_w_lg_reset_reconf_addr592w(0);
	wire_w_lg_w_lg_is_bonded_global_clk_div9w10w(0) <= wire_w_lg_is_bonded_global_clk_div9w(0) AND busy_state;
	wire_w_lg_w_lg_is_bonded_reconfig17w18w(0) <= wire_w_lg_is_bonded_reconfig17w(0) AND busy_state;
	wire_w_lg_w_lg_is_table_3313w14w(0) <= wire_w_lg_is_table_3313w(0) AND busy_state;
	wire_w_lg_w_lg_s2_to_058w59w(0) <= wire_w_lg_s2_to_058w(0) AND wire_w_lg_s0_to_157w(0);
	wire_w_lg_w_lg_s2_to_058w70w(0) <= wire_w_lg_s2_to_058w(0) AND wire_w_lg_s1_to_169w(0);
	wire_w_lg_w_lg_tx_reconfig93w94w(0) <= wire_w_lg_tx_reconfig93w(0) AND wire_w_lg_rx_reconfig92w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range842w850w851w(0) <= wire_w_lg_w_rx_eqctrl_range842w850w(0) AND wire_w_lg_w_rx_eqctrl_range840w841w(0);
	wire_w_lg_w_lg_w_w_rx_eqv959w_range1011w1018w1043w(0) <= wire_w_lg_w_w_rx_eqv959w_range1011w1018w(0) AND wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1041w1042w(0);
	wire_w_lg_w_lg_w_w_rx_eqv959w_range1011w1018w1054w(0) <= wire_w_lg_w_w_rx_eqv959w_range1011w1018w(0) AND wire_w_lg_w_w_rx_eqv959w_range1010w1017w(0);
	wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1019w1020w(0) <= wire_w_lg_w_w_rx_eqv959w_range1014w1019w(0) AND wire_w_lg_w_w_rx_eqv959w_range1011w1018w(0);
	wire_w_lg_w156w157w(0) <= wire_w156w(0) AND wire_w_lg_is_central_pcs149w(0);
	wire_w99w(0) <= wire_w_lg_w_lg_w_lg_w_lg_mif_type_error95w96w97w98w(0) AND write_state;
	loop5 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_w752w753w754w755w(i) <= wire_w_lg_w_lg_w752w753w754w(i) AND is_analog_control;
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_is_tier_1737w738w739w(i) <= wire_w_lg_w_lg_is_tier_1737w738w(0) AND reconfig_datain(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_dprio_datain_68_6B742w743w(i) <= wire_w_lg_dprio_datain_68_6B742w(i) AND write_word_68_6B_data_valid;
	END GENERATE loop7;
	wire_w_lg_w_lg_mif_type_error95w96w(0) <= wire_w_lg_mif_type_error95w(0) AND is_tier_1;
	wire_w_lg_w_lg_w_channel_address_range153w154w155w(0) <= wire_w_lg_w_channel_address_range153w154w(0) AND wire_w_lg_is_pll_address142w(0);
	wire_w_lg_w_lg_w_channel_address_range143w144w145w(0) <= wire_w_lg_w_channel_address_range143w144w(0) AND wire_w_lg_is_pll_address142w(0);
	wire_w_lg_w_lg_w_logical_pll_sel_num_range150w151w152w(0) <= wire_w_lg_w_logical_pll_sel_num_range150w151w(0) AND is_pll_address;
	wire_w_lg_w_lg_w_logical_pll_sel_num_range139w140w141w(0) <= wire_w_lg_w_logical_pll_sel_num_range139w140w(0) AND is_pll_address;
	wire_w_lg_adce_busy_state444w(0) <= adce_busy_state AND wire_w_adce_quad_addr_s4_range443w(0);
	wire_w_lg_adce_busy_state458w(0) <= adce_busy_state AND wire_w_adce_quad_addr_s4_range457w(0);
	wire_w_lg_adce_busy_state470w(0) <= adce_busy_state AND wire_w_adce_quad_addr_s4_range469w(0);
	wire_w_lg_adce_busy_state482w(0) <= adce_busy_state AND wire_w_adce_quad_addr_s4_range481w(0);
	wire_w_lg_adce_busy_state494w(0) <= adce_busy_state AND wire_w_adce_quad_addr_s4_range493w(0);
	wire_w_lg_adce_busy_state506w(0) <= adce_busy_state AND wire_w_adce_quad_addr_s4_range505w(0);
	loop8 : FOR i IN 0 TO 11 GENERATE 
		wire_w_lg_cal_busy186w(i) <= cal_busy AND wire_w185w(i);
	END GENERATE loop8;
	wire_w_lg_cal_busy516w(0) <= cal_busy AND wire_w_cal_quad_address_range515w(0);
	wire_w_lg_cal_busy525w(0) <= cal_busy AND wire_w_cal_quad_address_range524w(0);
	wire_w_lg_cal_busy533w(0) <= cal_busy AND wire_w_cal_quad_address_range532w(0);
	wire_w_lg_cal_busy541w(0) <= cal_busy AND wire_w_cal_quad_address_range540w(0);
	wire_w_lg_cal_busy549w(0) <= cal_busy AND wire_w_cal_quad_address_range548w(0);
	wire_w_lg_cal_busy557w(0) <= cal_busy AND wire_w_cal_quad_address_range556w(0);
	loop9 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_ctrl_address357w(i) <= ctrl_address(i) AND wire_w_lg_is_do_dfe356w(0);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_ctrl_address365w(i) <= ctrl_address(i) AND wire_w_lg_is_do_eyemon364w(0);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_ctrl_writedata360w(i) <= ctrl_writedata(i) AND wire_w_lg_is_do_dfe356w(0);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_ctrl_writedata368w(i) <= ctrl_writedata(i) AND wire_w_lg_is_do_eyemon364w(0);
	END GENERATE loop12;
	wire_w_lg_dfe_busy436w(0) <= dfe_busy AND wire_w_dfe_quad_address_range435w(0);
	wire_w_lg_dfe_busy452w(0) <= dfe_busy AND wire_w_dfe_quad_address_range451w(0);
	wire_w_lg_dfe_busy464w(0) <= dfe_busy AND wire_w_dfe_quad_address_range463w(0);
	wire_w_lg_dfe_busy476w(0) <= dfe_busy AND wire_w_dfe_quad_address_range475w(0);
	wire_w_lg_dfe_busy488w(0) <= dfe_busy AND wire_w_dfe_quad_address_range487w(0);
	wire_w_lg_dfe_busy500w(0) <= dfe_busy AND wire_w_dfe_quad_address_range499w(0);
	loop13 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain735w(i) <= dprio_datain(i) AND wire_w_lg_header_proc593w(0);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_64_67744w(i) <= dprio_datain_64_67(i) AND write_word_64_67_data_valid;
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_7c_7f741w(i) <= dprio_datain_7c_7f(i) AND write_word_7c_7f_data_valid;
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_7c_7f_inv740w(i) <= dprio_datain_7c_7f_inv(i) AND write_word_7c_7f_inv_data_valid;
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_preemp1t747w(i) <= dprio_datain_preemp1t(i) AND wire_w_lg_w_lg_write_word_preemp1t_data_valid745w746w(0);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_vodctrl749w(i) <= dprio_datain_vodctrl(i) AND wire_w_lg_write_word_vodctrl_data_valid748w(0);
	END GENERATE loop18;
	wire_w_lg_dprio_pulse709w(0) <= dprio_pulse AND wire_read_addr_cntr_w_lg_w_q_range693w708w(0);
	wire_w_lg_dprio_pulse716w(0) <= dprio_pulse AND wire_read_addr_cntr_w_q_range693w(0);
	wire_w_lg_eyemon_busy440w(0) <= eyemon_busy AND wire_w_eyemon_quad_address_range439w(0);
	wire_w_lg_eyemon_busy455w(0) <= eyemon_busy AND wire_w_eyemon_quad_address_range454w(0);
	wire_w_lg_eyemon_busy467w(0) <= eyemon_busy AND wire_w_eyemon_quad_address_range466w(0);
	wire_w_lg_eyemon_busy479w(0) <= eyemon_busy AND wire_w_eyemon_quad_address_range478w(0);
	wire_w_lg_eyemon_busy491w(0) <= eyemon_busy AND wire_w_eyemon_quad_address_range490w(0);
	wire_w_lg_eyemon_busy503w(0) <= eyemon_busy AND wire_w_eyemon_quad_address_range502w(0);
	wire_w_lg_idle_state50w(0) <= idle_state AND wire_w_lg_read49w(0);
	wire_w_lg_idle_state41w(0) <= idle_state AND wire_w_lg_w_lg_is_adce39w40w(0);
	loop19 : FOR i IN 0 TO 11 GENERATE 
		wire_w_lg_is_adce_mode_sel103w(i) <= is_adce_mode_sel AND default_max_limit_wire(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 11 GENERATE 
		wire_w_lg_is_analog_control108w(i) <= is_analog_control AND analog_write_max_limit(i);
	END GENERATE loop20;
	wire_w_lg_is_analog_control106w(0) <= is_analog_control AND read_state;
	wire_w_lg_is_bonded_reconfig23w(0) <= is_bonded_reconfig AND wire_w_lg_is_bonded_global_clk_div9w(0);
	wire_w_lg_is_bonded_reconfig16w(0) <= is_bonded_reconfig AND wire_w_lg_w_lg_w_lg_is_table_3313w14w15w(0);
	wire_w_lg_is_illegal_reg_d124w(0) <= is_illegal_reg_d AND wire_w_lg_w_lg_read_done120w123w(0);
	wire_w_lg_is_illegal_reg_out121w(0) <= is_illegal_reg_out AND wire_w_lg_read_done120w(0);
	wire_w_lg_is_table_3312w(0) <= is_table_33 AND wire_w_lg_w_lg_w_lg_is_bonded_global_clk_div9w10w11w(0);
	wire_w_lg_is_table_59138w(0) <= is_table_59 AND is_bonded_reconfig;
	wire_w_lg_is_table_61148w(0) <= is_table_61 AND is_central_pcs;
	wire_w_lg_is_tier_1613w(0) <= is_tier_1 AND wire_w_lg_header_proc593w(0);
	wire_w_lg_is_tier_1589w(0) <= is_tier_1 AND wire_w_lg_w587w588w(0);
	wire_w_lg_is_tier_1574w(0) <= is_tier_1 AND mif_reconfig_done;
	loop21 : FOR i IN 0 TO 11 GENERATE 
		wire_w_lg_is_tier_1105w(i) <= is_tier_1 AND tier_1_max_limit(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 11 GENERATE 
		wire_w_lg_is_tx_local_div_ctrl104w(i) <= is_tx_local_div_ctrl AND rate_switch_ctrl_max_limit(i);
	END GENERATE loop22;
	wire_w_lg_read49w(0) <= read AND en_read_trigger;
	loop23 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_read_address560w(i) <= read_address(i) AND read_state;
	END GENERATE loop23;
	wire_w_lg_read_state582w(0) <= read_state AND wire_w_lg_dprio_pulse581w(0);
	wire_w_lg_read_state1114w(0) <= read_state AND read_word_7c_7f_data_valid;
	loop24 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_read_state1068w(i) <= read_state AND w_rx_eqctrl_out954w(i);
	END GENERATE loop24;
	loop25 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_read_state1088w(i) <= read_state AND w_rx_eqdcgain_out1070w(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_read_state1111w(i) <= read_state AND w_tx_vodctrl_out1090w(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_read_state1124w(i) <= read_state AND wire_dprio_w_dataout_range797w(i);
	END GENERATE loop27;
	loop28 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_read_state1118w(i) <= read_state AND wire_dprio_w_dataout_range1117w(i);
	END GENERATE loop28;
	wire_w_lg_read_state1147w(0) <= read_state AND wire_dprio_w_dataout_range1146w(0);
	wire_w_lg_read_state1137w(0) <= read_state AND wire_dprio_w_dataout_range1136w(0);
	loop29 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_read_state1130w(i) <= read_state AND wire_dprio_w_dataout_range1129w(i);
	END GENERATE loop29;
	wire_w_lg_read_word_64_67_data_valid1085w(0) <= read_word_64_67_data_valid AND read_state;
	wire_w_lg_read_word_68_6B_data_valid1065w(0) <= read_word_68_6B_data_valid AND read_state;
	wire_w_lg_read_word_7c_7f_data_valid1126w(0) <= read_word_7c_7f_data_valid AND read_state;
	wire_w_lg_read_word_7c_7f_inv_data_valid703w(0) <= read_word_7c_7f_inv_data_valid AND wire_w_lg_rx_reconfig92w(0);
	wire_w_lg_read_word_preemp_1t_data_valid1121w(0) <= read_word_preemp_1t_data_valid AND read_state;
	wire_w_lg_read_word_vodctrl_data_valid1108w(0) <= read_word_vodctrl_data_valid AND read_state;
	loop30 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_eq_0_1004w1060w(i) <= w_eq_0_1004w(i) AND w_gt_0_only988w;
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_eq_10_1045w1057w(i) <= w_eq_10_1045w(i) AND w_gt_10_only1002w;
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_eq_3_1026w1059w(i) <= w_eq_3_1026w(i) AND w_gt_3_only995w;
	END GENERATE loop32;
	loop33 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_eq_6_1036w1058w(i) <= w_eq_6_1036w(i) AND w_gt_6_only999w;
	END GENERATE loop33;
	wire_w_lg_w_gt_0_964w992w(0) <= w_gt_0_964w AND wire_w_lg_w_gt_3_970w991w(0);
	wire_w_lg_w_gt_0_964w996w(0) <= w_gt_0_964w AND w_gt_3_970w;
	wire_w_lg_wr_pulse732w(0) <= wr_pulse AND wire_wren_data_reg_w_lg_q724w(0);
	wire_w_lg_wr_pulse729w(0) <= wr_pulse AND wire_wren_data_reg_w_lg_q728w(0);
	loop34 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_write_address561w(i) <= write_address(i) AND write_state;
	END GENERATE loop34;
	wire_w_lg_write_all25w(0) <= write_all AND wire_w_lg_w_lg_is_bonded_reconfig17w24w(0);
	wire_w_lg_write_state596w(0) <= write_state AND wire_w_lg_w_lg_w_lg_header_proc593w594w595w(0);
	wire_w_lg_write_state619w(0) <= write_state AND wire_w_lg_dprio_pulse581w(0);
	wire_w_lg_write_state1135w(0) <= write_state AND wire_w_lg_w_tx_preemp_0t_range2w896w(0);
	wire_w_lg_write_state1145w(0) <= write_state AND wire_w_lg_w_tx_preemp_2t_range4w900w(0);
	loop35 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_write_state1067w(i) <= write_state AND rx_eqctrl(i);
	END GENERATE loop35;
	loop36 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_write_state1087w(i) <= write_state AND rx_eqdcgain(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_write_state1123w(i) <= write_state AND tx_preemp_1t(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_write_state1110w(i) <= write_state AND tx_vodctrl(i);
	END GENERATE loop38;
	wire_w_lg_write_state1084w(0) <= write_state AND write_word_64_67_data_valid;
	wire_w_lg_write_state1064w(0) <= write_state AND write_word_68_6B_data_valid;
	wire_w_lg_write_state1113w(0) <= write_state AND write_word_7c_7f_data_valid;
	wire_w_lg_write_state1120w(0) <= write_state AND write_word_preemp1t_data_valid;
	wire_w_lg_write_state1107w(0) <= write_state AND write_word_vodctrl_data_valid;
	loop39 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_write_state1116w(i) <= write_state AND wire_w_tx_preemp_0t_wire_range894w(i);
	END GENERATE loop39;
	loop40 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_write_state1128w(i) <= write_state AND wire_w_tx_preemp_2t_wire_range898w(i);
	END GENERATE loop40;
	wire_w_lg_write_word_7c_7f_inv_data_valid938w(0) <= write_word_7c_7f_inv_data_valid AND wire_w_lg_rx_reconfig92w(0);
	wire_w_lg_write_word_done906w(0) <= write_word_done AND write_addr_inc;
	wire_w_lg_w_reconfig_mode_sel_range644w645w(0) <= wire_w_reconfig_mode_sel_range644w(0) AND wire_w_lg_w_reconfig_mode_sel_range85w643w(0);
	wire_w_lg_w_rx_eqctrl_range838w854w(0) <= wire_w_rx_eqctrl_range838w(0) AND wire_w_lg_w_rx_eqctrl_range845w853w(0);
	wire_w_lg_w_rx_eqctrl_range838w864w(0) <= wire_w_rx_eqctrl_range838w(0) AND wire_w_lg_w_rx_eqctrl_range845w863w(0);
	wire_w_lg_w_rx_eqctrl_range840w848w(0) <= wire_w_rx_eqctrl_range840w(0) AND wire_w_lg_w_rx_eqctrl_range838w839w(0);
	wire_w_lg_w_rx_eqctrl_range840w871w(0) <= wire_w_rx_eqctrl_range840w(0) AND wire_w_rx_eqctrl_range838w(0);
	wire_w_lg_w_rx_eqctrl_range842w843w(0) <= wire_w_rx_eqctrl_range842w(0) AND wire_w_lg_w_rx_eqctrl_range840w841w(0);
	wire_w_lg_w_rx_eqctrl_range842w869w(0) <= wire_w_rx_eqctrl_range842w(0) AND wire_w_rx_eqctrl_range838w(0);
	wire_w_lg_w_rx_eqctrl_range842w846w(0) <= wire_w_rx_eqctrl_range842w(0) AND wire_w_rx_eqctrl_range840w(0);
	wire_w_lg_w_rx_eqdcgain_range820w821w(0) <= wire_w_rx_eqdcgain_range820w(0) AND wire_w_rx_eqdcgain_range819w(0);
	wire_w_lg_w_tx_vodctrl_range761w769w(0) <= wire_w_tx_vodctrl_range761w(0) AND wire_w_lg_w_lg_w_tx_vodctrl_range759w760w768w(0);
	wire_w_lg_w_tx_vodctrl_range761w762w(0) <= wire_w_tx_vodctrl_range761w(0) AND wire_w_lg_w_tx_vodctrl_range759w760w(0);
	wire_w_lg_w_tx_vodctrl_range759w771w(0) <= wire_w_tx_vodctrl_range759w(0) AND wire_w_lg_w_tx_vodctrl_range758w770w(0);
	wire_w_lg_w_tx_vodctrl_range759w763w(0) <= wire_w_tx_vodctrl_range759w(0) AND wire_w_tx_vodctrl_range758w(0);
	wire_w_lg_w_w_rx_eqv959w_range1014w1015w(0) <= wire_w_w_rx_eqv959w_range1014w(0) AND wire_w_lg_w_lg_w_w_rx_eqv959w_range1011w1012w1013w(0);
	wire_w_lg_w_w_rx_eqv959w_range1014w1033w(0) <= wire_w_w_rx_eqv959w_range1014w(0) AND wire_w_lg_w_w_rx_eqv959w_range1011w1018w(0);
	wire_w_lg_w_w_rx_eqv959w_range1014w1022w(0) <= wire_w_w_rx_eqv959w_range1014w(0) AND wire_w_w_rx_eqv959w_range1011w(0);
	wire_w_lg_w_lg_read_done120w123w(0) <= NOT wire_w_lg_read_done120w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range842w873w874w(0) <= NOT wire_w_lg_w_rx_eqctrl_range842w873w(0);
	wire_w_lg_w_lg_w_tx_vodctrl_range759w760w768w(0) <= NOT wire_w_lg_w_tx_vodctrl_range759w760w(0);
	wire_w_lg_w_lg_w_w_rx_eqv959w_range1011w1012w1013w(0) <= NOT wire_w_lg_w_w_rx_eqv959w_range1011w1012w(0);
	wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1041w1042w(0) <= NOT wire_w_lg_w_w_rx_eqv959w_range1014w1041w(0);
	wire_w_lg_adce_busy_state132w(0) <= NOT adce_busy_state;
	wire_w_lg_bonded_skip604w(0) <= NOT bonded_skip;
	wire_w_lg_cal_busy182w(0) <= NOT cal_busy;
	wire_w_lg_dprio_pulse581w(0) <= NOT dprio_pulse;
	wire_w_lg_header_proc593w(0) <= NOT header_proc;
	wire_w_lg_idle_state117w(0) <= NOT idle_state;
	wire_w_lg_is_adce116w(0) <= NOT is_adce;
	wire_w_lg_is_analog_control731w(0) <= NOT is_analog_control;
	wire_w_lg_is_bonded_global_clk_div9w(0) <= NOT is_bonded_global_clk_div;
	wire_w_lg_is_bonded_reconfig17w(0) <= NOT is_bonded_reconfig;
	wire_w_lg_is_central_pcs149w(0) <= NOT is_central_pcs;
	wire_w_lg_is_cruclk_addr0606w(0) <= NOT is_cruclk_addr0;
	wire_w_lg_is_diff_mif564w(0) <= NOT is_diff_mif;
	wire_w_lg_is_do_dfe356w(0) <= NOT is_do_dfe;
	wire_w_lg_is_do_eyemon364w(0) <= NOT is_do_eyemon;
	wire_w_lg_is_global_clk_div_mode602w(0) <= NOT is_global_clk_div_mode;
	wire_w_lg_is_illegal_reg_d579w(0) <= NOT is_illegal_reg_d;
	wire_w_lg_is_illegal_reg_out122w(0) <= NOT is_illegal_reg_out;
	wire_w_lg_is_pll_address142w(0) <= NOT is_pll_address;
	wire_w_lg_is_protected_bit603w(0) <= NOT is_protected_bit;
	wire_w_lg_is_rcxpat_chnl_en_ch607w(0) <= NOT is_rcxpat_chnl_en_ch;
	wire_w_lg_is_table_3313w(0) <= NOT is_table_33;
	wire_w_lg_is_tier_1590w(0) <= NOT is_tier_1;
	wire_w_lg_rd_pulse198w(0) <= NOT rd_pulse;
	wire_w_lg_read_done580w(0) <= NOT read_done;
	wire_w_lg_read_state571w(0) <= NOT read_state;
	wire_w_lg_reconfig_reset_all28w(0) <= NOT reconfig_reset_all;
	wire_w_lg_reset_reconf_addr592w(0) <= NOT reset_reconf_addr;
	wire_w_lg_rx_reconfig92w(0) <= NOT rx_reconfig;
	wire_w_lg_s0_to_056w(0) <= NOT s0_to_0;
	wire_w_lg_s0_to_157w(0) <= NOT s0_to_1;
	wire_w_lg_s1_to_068w(0) <= NOT s1_to_0;
	wire_w_lg_s1_to_169w(0) <= NOT s1_to_1;
	wire_w_lg_s2_to_058w(0) <= NOT s2_to_0;
	wire_w_lg_tx_reconfig93w(0) <= NOT tx_reconfig;
	wire_w_lg_w_gt_10_982w989w(0) <= NOT w_gt_10_982w;
	wire_w_lg_w_gt_3_970w991w(0) <= NOT w_gt_3_970w;
	wire_w_lg_w_gt_6_976w990w(0) <= NOT w_gt_6_976w;
	wire_w_lg_wr_pulse199w(0) <= NOT wr_pulse;
	wire_w_lg_write_all_int47w(0) <= NOT write_all_int;
	wire_w_lg_write_done91w(0) <= NOT write_done;
	wire_w_lg_write_skip605w(0) <= NOT write_skip;
	wire_w_lg_write_state48w(0) <= NOT write_state;
	wire_w_lg_w_reconfig_mode_sel_range85w643w(0) <= NOT wire_w_reconfig_mode_sel_range85w(0);
	wire_w_lg_w_rx_eqctrl_range845w853w(0) <= NOT wire_w_rx_eqctrl_range845w(0);
	wire_w_lg_w_rx_eqctrl_range838w839w(0) <= NOT wire_w_rx_eqctrl_range838w(0);
	wire_w_lg_w_rx_eqctrl_range840w841w(0) <= NOT wire_w_rx_eqctrl_range840w(0);
	wire_w_lg_w_rx_eqctrl_range842w850w(0) <= NOT wire_w_rx_eqctrl_range842w(0);
	wire_w_lg_w_tx_preemp_0t_range2w896w(0) <= NOT wire_w_tx_preemp_0t_range2w(0);
	wire_w_lg_w_tx_preemp_2t_range4w900w(0) <= NOT wire_w_tx_preemp_2t_range4w(0);
	wire_w_lg_w_tx_vodctrl_range758w770w(0) <= NOT wire_w_tx_vodctrl_range758w(0);
	wire_w_lg_w_w_rx_eqv959w_range1010w1017w(0) <= NOT wire_w_w_rx_eqv959w_range1010w(0);
	wire_w_lg_w_w_rx_eqv959w_range1011w1018w(0) <= NOT wire_w_w_rx_eqv959w_range1011w(0);
	wire_w_lg_w_w_rx_eqv959w_range1014w1019w(0) <= NOT wire_w_w_rx_eqv959w_range1014w(0);
	wire_w_lg_w876w877w(0) <= wire_w876w(0) OR wire_w_lg_w_lg_w_rx_eqctrl_range840w871w872w(0);
	wire_w1024w(0) <= wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1022w1023w(0) OR wire_w1021w(0);
	wire_w_lg_w_lg_w_lg_cal_busy182w511w512w(0) <= wire_w_lg_w_lg_cal_busy182w511w(0) OR wire_w_w_wire_eyemon_dprioout_mux432w_range441w(0);
	wire_w_lg_w_lg_w_lg_cal_busy182w520w521w(0) <= wire_w_lg_w_lg_cal_busy182w520w(0) OR wire_w_w_wire_eyemon_dprioout_mux432w_range456w(0);
	wire_w_lg_w_lg_w_lg_cal_busy182w528w529w(0) <= wire_w_lg_w_lg_cal_busy182w528w(0) OR wire_w_w_wire_eyemon_dprioout_mux432w_range468w(0);
	wire_w_lg_w_lg_w_lg_cal_busy182w536w537w(0) <= wire_w_lg_w_lg_cal_busy182w536w(0) OR wire_w_w_wire_eyemon_dprioout_mux432w_range480w(0);
	wire_w_lg_w_lg_w_lg_cal_busy182w544w545w(0) <= wire_w_lg_w_lg_cal_busy182w544w(0) OR wire_w_w_wire_eyemon_dprioout_mux432w_range492w(0);
	wire_w_lg_w_lg_w_lg_cal_busy182w552w553w(0) <= wire_w_lg_w_lg_cal_busy182w552w(0) OR wire_w_w_wire_eyemon_dprioout_mux432w_range504w(0);
	wire_w_lg_w_lg_w_lg_is_bonded_global_clk_div9w10w11w(0) <= wire_w_lg_w_lg_is_bonded_global_clk_div9w10w(0) OR is_bonded_global_clk_div;
	wire_w_lg_w_lg_w_lg_is_table_3313w14w15w(0) <= wire_w_lg_w_lg_is_table_3313w14w(0) OR wire_w_lg_is_table_3312w(0);
	wire_w1052w(0) <= wire_w_lg_w_lg_w_w_rx_eqv959w_range1011w1018w1043w(0) OR wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1022w1023w(0);
	wire_w1055w(0) <= wire_w_lg_w_lg_w_w_rx_eqv959w_range1011w1018w1054w(0) OR wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1022w1023w(0);
	wire_w_lg_w_lg_w156w157w158w(0) <= wire_w_lg_w156w157w(0) OR wire_w_lg_is_table_61148w(0);
	wire_w_lg_w_lg_w_lg_mif_type_error95w96w97w(0) <= wire_w_lg_w_lg_mif_type_error95w96w(0) OR wire_w_lg_w_lg_tx_reconfig93w94w(0);
	wire_w156w(0) <= wire_w_lg_w_lg_w_channel_address_range153w154w155w(0) OR wire_w_lg_w_lg_w_logical_pll_sel_num_range150w151w152w(0);
	wire_w146w(0) <= wire_w_lg_w_lg_w_channel_address_range143w144w145w(0) OR wire_w_lg_w_lg_w_logical_pll_sel_num_range139w140w141w(0);
	loop41 : FOR i IN 0 TO 11 GENERATE 
		wire_w_lg_w_lg_cal_busy186w187w(i) <= wire_w_lg_cal_busy186w(i) OR wire_w_lg_w_lg_cal_busy182w183w(i);
	END GENERATE loop41;
	wire_w_lg_w_lg_cal_busy516w517w(0) <= wire_w_lg_cal_busy516w(0) OR wire_w514w(0);
	wire_w_lg_w_lg_cal_busy525w526w(0) <= wire_w_lg_cal_busy525w(0) OR wire_w523w(0);
	wire_w_lg_w_lg_cal_busy533w534w(0) <= wire_w_lg_cal_busy533w(0) OR wire_w531w(0);
	wire_w_lg_w_lg_cal_busy541w542w(0) <= wire_w_lg_cal_busy541w(0) OR wire_w539w(0);
	wire_w_lg_w_lg_cal_busy549w550w(0) <= wire_w_lg_cal_busy549w(0) OR wire_w547w(0);
	wire_w_lg_w_lg_cal_busy557w558w(0) <= wire_w_lg_cal_busy557w(0) OR wire_w555w(0);
	loop42 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_dprio_datain_vodctrl749w750w(i) <= wire_w_lg_dprio_datain_vodctrl749w(i) OR wire_w_lg_dprio_datain_preemp1t747w(i);
	END GENERATE loop42;
	wire_w_lg_w_lg_read_state1114w1115w(0) <= wire_w_lg_read_state1114w(0) OR wire_w_lg_write_state1113w(0);
	loop43 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_lg_read_state1068w1069w(i) <= wire_w_lg_read_state1068w(i) OR wire_w_lg_write_state1067w(i);
	END GENERATE loop43;
	loop44 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_w_lg_read_state1088w1089w(i) <= wire_w_lg_read_state1088w(i) OR wire_w_lg_write_state1087w(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 2 GENERATE 
		wire_w_lg_w_lg_read_state1111w1112w(i) <= wire_w_lg_read_state1111w(i) OR wire_w_lg_write_state1110w(i);
	END GENERATE loop45;
	loop46 : FOR i IN 0 TO 4 GENERATE 
		wire_w_lg_w_lg_read_state1124w1125w(i) <= wire_w_lg_read_state1124w(i) OR wire_w_lg_write_state1123w(i);
	END GENERATE loop46;
	loop47 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_lg_read_state1118w1119w(i) <= wire_w_lg_read_state1118w(i) OR wire_w_lg_write_state1116w(i);
	END GENERATE loop47;
	loop48 : FOR i IN 0 TO 3 GENERATE 
		wire_w_lg_w_lg_read_state1130w1131w(i) <= wire_w_lg_read_state1130w(i) OR wire_w_lg_write_state1128w(i);
	END GENERATE loop48;
	wire_w_lg_w_lg_read_word_64_67_data_valid1085w1086w(0) <= wire_w_lg_read_word_64_67_data_valid1085w(0) OR wire_w_lg_write_state1084w(0);
	wire_w_lg_w_lg_read_word_68_6B_data_valid1065w1066w(0) <= wire_w_lg_read_word_68_6B_data_valid1065w(0) OR wire_w_lg_write_state1064w(0);
	wire_w_lg_w_lg_read_word_7c_7f_data_valid1126w1127w(0) <= wire_w_lg_read_word_7c_7f_data_valid1126w(0) OR wire_w_lg_write_state1113w(0);
	wire_w_lg_w_lg_read_word_preemp_1t_data_valid1121w1122w(0) <= wire_w_lg_read_word_preemp_1t_data_valid1121w(0) OR wire_w_lg_write_state1120w(0);
	wire_w_lg_w_lg_read_word_vodctrl_data_valid1108w1109w(0) <= wire_w_lg_read_word_vodctrl_data_valid1108w(0) OR wire_w_lg_write_state1107w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range838w854w855w(0) <= wire_w_lg_w_rx_eqctrl_range838w854w(0) OR wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range842w850w851w852w(0);
	wire_w_lg_w_lg_w_rx_eqctrl_range838w864w865w(0) <= wire_w_lg_w_rx_eqctrl_range838w864w(0) OR wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range842w846w860w861w(0);
	wire_w_lg_w_lg_w_tx_vodctrl_range759w771w772w(0) <= wire_w_lg_w_tx_vodctrl_range759w771w(0) OR wire_w_lg_w_tx_vodctrl_range761w769w(0);
	wire_w_lg_w_lg_w_tx_vodctrl_range759w763w764w(0) <= wire_w_lg_w_tx_vodctrl_range759w763w(0) OR wire_w_lg_w_tx_vodctrl_range761w762w(0);
	wire_w_lg_w_lg_is_bonded_reconfig17w24w(0) <= wire_w_lg_is_bonded_reconfig17w(0) OR wire_w_lg_is_bonded_reconfig23w(0);
	wire_w_lg_w_lg_is_tier_1590w616w(0) <= wire_w_lg_is_tier_1590w(0) OR wire_w_lg_w_lg_is_tier_1613w615w(0);
	wire_w_lg_w_lg_is_tier_1590w591w(0) <= wire_w_lg_is_tier_1590w(0) OR wire_w_lg_is_tier_1589w(0);
	wire_w_lg_w_lg_w876w877w878w(0) <= wire_w_lg_w876w877w(0) OR wire_w_lg_w_lg_w_rx_eqctrl_range842w869w870w(0);
	wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w511w512w513w(0) <= wire_w_lg_w_lg_w_lg_cal_busy182w511w512w(0) OR wire_w_w_wire_adce_dprioout_mux433w_range445w(0);
	wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w520w521w522w(0) <= wire_w_lg_w_lg_w_lg_cal_busy182w520w521w(0) OR wire_w_w_wire_adce_dprioout_mux433w_range459w(0);
	wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w528w529w530w(0) <= wire_w_lg_w_lg_w_lg_cal_busy182w528w529w(0) OR wire_w_w_wire_adce_dprioout_mux433w_range471w(0);
	wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w536w537w538w(0) <= wire_w_lg_w_lg_w_lg_cal_busy182w536w537w(0) OR wire_w_w_wire_adce_dprioout_mux433w_range483w(0);
	wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w544w545w546w(0) <= wire_w_lg_w_lg_w_lg_cal_busy182w544w545w(0) OR wire_w_w_wire_adce_dprioout_mux433w_range495w(0);
	wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w552w553w554w(0) <= wire_w_lg_w_lg_w_lg_cal_busy182w552w553w(0) OR wire_w_w_wire_adce_dprioout_mux433w_range507w(0);
	wire_w_lg_w_lg_w_lg_w_lg_mif_type_error95w96w97w98w(0) <= wire_w_lg_w_lg_w_lg_mif_type_error95w96w97w(0) OR invalid_eq_dcgain;
	wire_w_lg_w146w147w(0) <= wire_w146w(0) OR is_central_pcs;
	loop49 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w_lg_dprio_datain_vodctrl749w750w751w(i) <= wire_w_lg_w_lg_dprio_datain_vodctrl749w750w(i) OR wire_w_lg_dprio_datain_64_67744w(i);
	END GENERATE loop49;
	wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range838w854w855w856w(0) <= wire_w_lg_w_lg_w_rx_eqctrl_range838w854w855w(0) OR wire_w_lg_w_lg_w_rx_eqctrl_range840w848w849w(0);
	wire_w_lg_w_lg_w_lg_w876w877w878w879w(0) <= wire_w_lg_w_lg_w876w877w878w(0) OR wire_w_lg_w_lg_w_rx_eqctrl_range842w846w868w(0);
	wire_w514w(0) <= wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w511w512w513w(0) OR wire_w_w_wire_adce_dprioout_mux2434w_range449w(0);
	wire_w523w(0) <= wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w520w521w522w(0) OR wire_w_w_wire_adce_dprioout_mux2434w_range462w(0);
	wire_w531w(0) <= wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w528w529w530w(0) OR wire_w_w_wire_adce_dprioout_mux2434w_range474w(0);
	wire_w539w(0) <= wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w536w537w538w(0) OR wire_w_w_wire_adce_dprioout_mux2434w_range486w(0);
	wire_w547w(0) <= wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w544w545w546w(0) OR wire_w_w_wire_adce_dprioout_mux2434w_range498w(0);
	wire_w555w(0) <= wire_w_lg_w_lg_w_lg_w_lg_cal_busy182w552w553w554w(0) OR wire_w_w_wire_adce_dprioout_mux2434w_range510w(0);
	loop50 : FOR i IN 0 TO 15 GENERATE 
		wire_w752w(i) <= wire_w_lg_w_lg_w_lg_dprio_datain_vodctrl749w750w751w(i) OR wire_w_lg_w_lg_dprio_datain_68_6B742w743w(i);
	END GENERATE loop50;
	wire_w857w(0) <= wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range838w854w855w856w(0) OR wire_w_lg_w_lg_w_rx_eqctrl_range842w846w847w(0);
	wire_w_lg_w_lg_w_lg_w_lg_w876w877w878w879w880w(0) <= wire_w_lg_w_lg_w_lg_w876w877w878w879w(0) OR wire_w_lg_w_lg_w_lg_w_rx_eqctrl_range842w843w844w867w(0);
	loop51 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w752w753w(i) <= wire_w752w(i) OR wire_w_lg_dprio_datain_7c_7f741w(i);
	END GENERATE loop51;
	wire_w_lg_w857w858w(0) <= wire_w857w(0) OR wire_w_lg_w_lg_w_rx_eqctrl_range842w843w844w(0);
	loop52 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_w_lg_w752w753w754w(i) <= wire_w_lg_w752w753w(i) OR wire_w_lg_dprio_datain_7c_7f_inv740w(i);
	END GENERATE loop52;
	wire_w_lg_w587w588w(0) <= wire_w587w(0) OR is_global_clk_div_mode;
	wire_w587w(0) <= wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch584w585w586w(0) OR is_protected_bit;
	wire_w_lg_w_lg_w_lg_is_rcxpat_chnl_en_ch584w585w586w(0) <= wire_w_lg_w_lg_is_rcxpat_chnl_en_ch584w585w(0) OR bonded_skip;
	wire_w_lg_w_lg_is_adce39w40w(0) <= wire_w_lg_is_adce39w(0) OR is_do_dfe;
	wire_w_lg_w_lg_is_pll_address135w136w(0) <= wire_w_lg_is_pll_address135w(0) OR is_bonded_global_clk_div;
	wire_w_lg_w_lg_is_rcxpat_chnl_en_ch584w585w(0) <= wire_w_lg_is_rcxpat_chnl_en_ch584w(0) OR write_skip;
	wire_w_lg_w_lg_is_tier_1737w738w(0) <= wire_w_lg_is_tier_1737w(0) OR is_tx_local_div_ctrl;
	wire_w_lg_w_lg_s0_to_262w63w(0) <= wire_w_lg_s0_to_262w(0) OR wire_w_lg_w_lg_w_lg_w_lg_s2_to_058w59w60w61w(0);
	wire_w_lg_w_lg_s0_to_273w74w(0) <= wire_w_lg_s0_to_273w(0) OR wire_w_lg_w_lg_w_lg_w_lg_s2_to_058w70w71w72w(0);
	wire_w_lg_w_lg_write_word_preemp1t_data_valid745w746w(0) <= wire_w_lg_write_word_preemp1t_data_valid745w(0) OR write_word_preemp1tb_data_valid;
	wire_w_lg_w_lg_w_rx_eqdcgain_range816w824w826w(0) <= wire_w_lg_w_rx_eqdcgain_range816w824w(0) OR wire_w_rx_eqdcgain_range819w(0);
	wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1049w1050w(0) <= wire_w_lg_w_w_rx_eqv959w_range1014w1049w(0) OR wire_w_w_rx_eqv959w_range1010w(0);
	wire_w_lg_adce_busy_state128w(0) <= adce_busy_state OR is_do_eyemon;
	loop53 : FOR i IN 0 TO 15 GENERATE 
		wire_w_lg_dprio_datain_68_6B742w(i) <= dprio_datain_68_6B(i) OR local_ch_dec;
	END GENERATE loop53;
	wire_w_lg_is_adce39w(0) <= is_adce OR is_do_eyemon;
	wire_w_lg_is_do_eyemon131w(0) <= is_do_eyemon OR is_do_dfe;
	wire_w_lg_is_pll_address135w(0) <= is_pll_address OR is_central_pcs;
	wire_w_lg_is_rcxpat_chnl_en_ch584w(0) <= is_rcxpat_chnl_en_ch OR is_cruclk_addr0;
	wire_w_lg_is_tier_1737w(0) <= is_tier_1 OR is_tier_2;
	wire_w_lg_mif_type_error95w(0) <= mif_type_error OR mif_family_error;
	wire_w_lg_read_done120w(0) <= read_done OR write_done;
	wire_w_lg_reset_system575w(0) <= reset_system OR wire_w_lg_is_tier_1574w(0);
	wire_w_lg_s0_to_262w(0) <= s0_to_2 OR s0_to_1;
	wire_w_lg_s0_to_273w(0) <= s0_to_2 OR s1_to_1;
	wire_w_lg_write_word_preemp1t_data_valid745w(0) <= write_word_preemp1t_data_valid OR write_word_preemp1ta_data_valid;
	wire_w_lg_write_word_vodctrl_data_valid748w(0) <= write_word_vodctrl_data_valid OR write_word_vodctrla_data_valid;
	wire_w_lg_w_channel_address_range153w154w(0) <= wire_w_channel_address_range153w(0) OR is_bonded_global_clk_div;
	wire_w_lg_w_channel_address_range143w144w(0) <= wire_w_channel_address_range143w(0) OR is_bonded_global_clk_div;
	wire_w_lg_w_logical_pll_sel_num_range150w151w(0) <= wire_w_logical_pll_sel_num_range150w(0) OR wire_w_lg_is_table_59138w(0);
	wire_w_lg_w_logical_pll_sel_num_range139w140w(0) <= wire_w_logical_pll_sel_num_range139w(0) OR wire_w_lg_is_table_59138w(0);
	wire_w_lg_w_rx_eqdcgain_range816w822w(0) <= wire_w_rx_eqdcgain_range816w(0) OR wire_w_lg_w_rx_eqdcgain_range820w821w(0);
	wire_w_lg_w_rx_eqdcgain_range816w824w(0) <= wire_w_rx_eqdcgain_range816w(0) OR wire_w_rx_eqdcgain_range820w(0);
	wire_w_lg_w_w_rx_eqv959w_range1014w1049w(0) <= wire_w_w_rx_eqv959w_range1014w(0) OR wire_w_w_rx_eqv959w_range1011w(0);
	wire_w_lg_w_rx_eqctrl_range845w863w(0) <= wire_w_rx_eqctrl_range845w(0) XOR wire_w_lg_w_rx_eqctrl_range840w862w(0);
	wire_w_lg_w_rx_eqctrl_range840w862w(0) <= wire_w_rx_eqctrl_range840w(0) XOR wire_w_rx_eqctrl_range842w(0);
	wire_w_lg_w_rx_eqctrl_range842w873w(0) <= wire_w_rx_eqctrl_range842w(0) XOR wire_w_rx_eqctrl_range840w(0);
	wire_w_lg_w_tx_vodctrl_range759w760w(0) <= wire_w_tx_vodctrl_range759w(0) XOR wire_w_tx_vodctrl_range758w(0);
	wire_w_lg_w_w_rx_eqv959w_range1011w1012w(0) <= wire_w_w_rx_eqv959w_range1011w(0) XOR wire_w_w_rx_eqv959w_range1010w(0);
	wire_w_lg_w_w_rx_eqv959w_range1014w1041w(0) <= wire_w_w_rx_eqv959w_range1014w(0) XOR wire_w_w_rx_eqv959w_range1010w(0);
	a2gr_dprio_addr <= (wire_w_lg_write_address561w OR wire_w_lg_read_address560w);
	a2gr_dprio_data <= wire_w_lg_w_lg_dprio_datain735w736w;
	a2gr_dprio_rden <= (rd_pulse AND (wire_w_lg_is_diff_mif564w(0) OR (is_diff_mif AND diff_mif_wr_rd_busy)));
	a2gr_dprio_wren <= ((wire_w_lg_wr_pulse732w(0) AND wire_w_lg_is_analog_control731w(0)) AND (wire_w_lg_is_diff_mif564w(0) OR (is_diff_mif AND diff_mif_wr_rd_busy)));
	a2gr_dprio_wren_data <= (wire_w_lg_wr_pulse729w(0) AND (wire_w_lg_is_diff_mif564w(0) OR (is_diff_mif AND diff_mif_wr_rd_busy)));
	adce_busy_state <= '0';
	adce_error_wire <= '0';
	adce_pres_reg <= (OTHERS => '0');
	adce_quad_addr_s4 <= (OTHERS => '0');
	adce_state <= (state_mc_reg(0) AND state_mc_reg(1));
	aeq_ch_done <= (OTHERS => '0');
	analog_read_max_limit <= "011011000000";
	analog_write_max_limit <= "110110000000";
	bonded_skip <= '0';
	busy <= (((wire_w_lg_w_lg_is_bonded_reconfig17w18w(0) OR wire_w_lg_is_bonded_reconfig16w(0)) OR internal_write_pulse) OR cal_busy);
	busy_state <= ((((read_state OR write_state) OR adce_state) OR eyemon_busy) OR dfe_busy);
	cal_busy <= wire_calibration_busy;
	cal_channel_address <= wire_calibration_dprio_addr(14 DOWNTO 12);
	cal_channel_address_out <= address_pres_reg(2 DOWNTO 0);
	cal_dprio_address <= ( wire_calibration_dprio_addr(15) & cal_channel_address_out & wire_calibration_dprio_addr(11 DOWNTO 0));
	cal_dprioout_wire <= ( reconfig_fromgxb(595) & reconfig_fromgxb(578) & reconfig_fromgxb(561) & reconfig_fromgxb(544) & reconfig_fromgxb(527) & reconfig_fromgxb(510) & reconfig_fromgxb(493) & reconfig_fromgxb(476) & reconfig_fromgxb(459) & reconfig_fromgxb(442) & reconfig_fromgxb(425) & reconfig_fromgxb(408) & reconfig_fromgxb(391) & reconfig_fromgxb(374) & reconfig_fromgxb(357) & reconfig_fromgxb(340) & reconfig_fromgxb(323) & reconfig_fromgxb(306) & reconfig_fromgxb(289) & reconfig_fromgxb(272) & reconfig_fromgxb(255) & reconfig_fromgxb(238) & reconfig_fromgxb(221) & reconfig_fromgxb(204) & reconfig_fromgxb(187) & reconfig_fromgxb(170) & reconfig_fromgxb(153) & reconfig_fromgxb(136) & reconfig_fromgxb(119) & reconfig_fromgxb(102) & reconfig_fromgxb(85) & reconfig_fromgxb(68) & reconfig_fromgxb(51) & reconfig_fromgxb(34) & reconfig_fromgxb(17) & reconfig_fromgxb(0));
	cal_quad_address <= wire_calibration_quad_addr;
	cal_testbuses <= ( reconfig_fromgxb(611 DOWNTO 596) & reconfig_fromgxb(594 DOWNTO 579) & reconfig_fromgxb(577 DOWNTO 562) & reconfig_fromgxb(560 DOWNTO 545) & reconfig_fromgxb(543 DOWNTO 528) & reconfig_fromgxb(526 DOWNTO 511) & reconfig_fromgxb(509 DOWNTO 494) & reconfig_fromgxb(492 DOWNTO 477) & reconfig_fromgxb(475 DOWNTO 460) & reconfig_fromgxb(458 DOWNTO 443) & reconfig_fromgxb(441 DOWNTO 426) & reconfig_fromgxb(424 DOWNTO 409) & reconfig_fromgxb(407 DOWNTO 392) & reconfig_fromgxb(390 DOWNTO 375) & reconfig_fromgxb(373 DOWNTO 358) & reconfig_fromgxb(356 DOWNTO 341) & reconfig_fromgxb(339 DOWNTO 324) & reconfig_fromgxb(322 DOWNTO 307) & reconfig_fromgxb(305 DOWNTO 290) & reconfig_fromgxb(288 DOWNTO 273) & reconfig_fromgxb(271 DOWNTO 256) & reconfig_fromgxb(254 DOWNTO 239) & reconfig_fromgxb(237 DOWNTO 222) & reconfig_fromgxb(220 DOWNTO 205) & reconfig_fromgxb(203 DOWNTO 188) & reconfig_fromgxb(186 DOWNTO 171) & reconfig_fromgxb(169 DOWNTO 154) & reconfig_fromgxb(152 DOWNTO 137) & reconfig_fromgxb(135 DOWNTO 120) & reconfig_fromgxb(118 DOWNTO 103) & reconfig_fromgxb(101 DOWNTO 86) & reconfig_fromgxb(84 DOWNTO 69) & reconfig_fromgxb(67 DOWNTO 52) & reconfig_fromgxb(50 DOWNTO 35) & reconfig_fromgxb(33 DOWNTO 18) & reconfig_fromgxb(16 DOWNTO 1));
	channel_address <= wire_addr_cntr_q(1 DOWNTO 0);
	channel_address_out <= wire_address_pres_reg_w_lg_w_q_range195w196w;
	ctrl_readdata <= (eyemon_readdata OR dfe_readdata);
	ctrl_waitrequest <= (eyemon_swaitrequest OR dfe_swaitrequest);
	data_valid <= (data_valid_reg AND idle_state);
	default_max_limit_wire <= "011111100000";
	dfe_busy <= wire_dfe_o_reconfig_busy;
	dfe_dprio_addr <= wire_dfe_o_dprio_addr;
	dfe_dprio_data <= wire_dfe_o_dprio_data;
	dfe_dprio_rden <= wire_dfe_o_dprio_rden;
	dfe_dprio_wren <= wire_dfe_o_dprio_wren;
	dfe_pres_reg <= ( wire_dfe_o_quad_address & "0" & wire_dfe_o_dprio_addr(13 DOWNTO 12));
	dfe_quad_address <= wire_dfe_o_quad_address;
	dfe_readdata <= wire_dfe_o_avmm_sreaddata;
	dfe_swaitrequest <= wire_dfe_o_avmm_swaitrequest;
	diff_mif_wr_rd_busy <= '0';
	dprio_datain <= (wire_w_lg_w_lg_w_lg_w752w753w754w755w OR wire_w_lg_w_lg_w_lg_is_tier_1737w738w739w);
	dprio_datain_64_67 <= ( wire_dprio_dataout(15 DOWNTO 11) & ( rx_eqdcgain(2) & wire_w_lg_w_rx_eqdcgain_range816w822w & wire_w_lg_w_rx_eqdcgain_range816w824w & wire_w_lg_w_lg_w_rx_eqdcgain_range816w824w826w) & wire_dprio_dataout(6 DOWNTO 0));
	dprio_datain_68_6B <= ( wire_dprio_dataout(15) & ( wire_cmpr7_agb & wire_cmpr7_agb & wire_cmpr7_agb & wire_cmpr8_agb & wire_cmpr8_agb & wire_cmpr8_agb & wire_cmpr9_agb & wire_cmpr9_agb & wire_cmpr9_agb & wire_cmpr10_agb & wire_cmpr10_agb & wire_cmpr10_agb & wire_w_lg_w857w858w & wire_w_lg_w_lg_w_rx_eqctrl_range838w864w865w & wire_w_lg_w_lg_w_lg_w_lg_w876w877w878w879w880w));
	dprio_datain_7c_7f <= ( wire_dprio_dataout(15 DOWNTO 8) & tx_preemp_2t_wire(3 DOWNTO 0) & tx_preemp_0t_wire(3 DOWNTO 0));
	dprio_datain_7c_7f_inv <= ( wire_dprio_dataout(15 DOWNTO 5) & wire_w_lg_w_tx_preemp_0t_range2w896w & wire_w_lg_w_tx_preemp_2t_range4w900w & wire_dprio_dataout(2 DOWNTO 0));
	dprio_datain_preemp1t <= ( tx_preemp_1t & wire_dprio_dataout(10 DOWNTO 0));
	dprio_datain_vodctrl <= ( ( wire_w_lg_w_lg_w_tx_vodctrl_range759w763w764w & wire_w_lg_w_tx_vodctrl_range759w760w & wire_w_lg_w_lg_w_tx_vodctrl_range759w771w772w) & wire_dprio_dataout(12 DOWNTO 0));
	dprio_pulse <= ((dprio_pulse_reg XOR wire_dprio_busy) AND wire_dprio_w_lg_busy567w(0));
	en_read_trigger <= '1';
	en_write_trigger <= '1';
	error <= error_reg;
	eyemon_busy <= wire_eyemonitor_o_reconfig_busy;
	eyemon_dprio_addr <= wire_eyemonitor_o_dprio_addr;
	eyemon_dprio_data <= wire_eyemonitor_o_dprio_data;
	eyemon_dprio_rden <= wire_eyemonitor_o_dprio_rden;
	eyemon_dprio_wren <= wire_eyemonitor_o_dprio_wren;
	eyemon_pres_reg <= ( wire_eyemonitor_o_quad_address & wire_eyemonitor_o_dprio_addr(14 DOWNTO 12));
	eyemon_quad_address <= wire_eyemonitor_o_quad_address;
	eyemon_readdata <= wire_eyemonitor_o_avmm_sreaddata;
	eyemon_swaitrequest <= wire_eyemonitor_o_avmm_swaitrequest;
	header_proc <= '0';
	idle_state <= (wire_state_mc_reg_w_lg_q31w(0) AND wire_state_mc_reg_w_lg_q29w(0));
	internal_write_pulse <= '0';
	invalid_eq_dcgain <= '0';
	is_adce <= ((((is_adce_single_control OR is_adce_all_control) OR is_adce_continuous_single_control) OR is_adce_one_time_single_control) OR is_adce_standby_single_control);
	is_adce_all_control <= '0';
	is_adce_continuous_single_control <= '0';
	is_adce_mode_sel <= ((wire_reconf_mode_dec_eq(8) OR wire_reconf_mode_dec_eq(9)) OR wire_reconf_mode_dec_eq(10));
	is_adce_one_time_single_control <= '0';
	is_adce_single_control <= '0';
	is_adce_standby_single_control <= '0';
	is_analog_control <= wire_reconf_mode_dec_eq(0);
	is_bonded_global_clk_div <= '0';
	is_bonded_reconfig <= '0';
	is_central_pcs <= '0';
	is_cruclk_addr0 <= '0';
	is_diff_mif <= '0';
	is_do_dfe <= ((((NOT reconfig_mode_sel(0)) AND wire_w_lg_w_reconfig_mode_sel_range85w643w(0)) AND reconfig_mode_sel(2)) AND reconfig_mode_sel(3));
	is_do_eyemon <= ((((reconfig_mode_sel(0) AND reconfig_mode_sel(1)) AND (NOT reconfig_mode_sel(2))) AND reconfig_mode_sel(3)) OR ((wire_w_lg_w_reconfig_mode_sel_range644w645w(0) AND reconfig_mode_sel(2)) AND reconfig_mode_sel(3)));
	is_global_clk_div_mode <= '0';
	is_illegal_reg_d <= ((((((is_tier_2 OR is_adce_mode_sel) OR (is_tier_1 AND read_state)) OR (is_tx_local_div_ctrl AND write_state)) OR (is_tx_local_div_ctrl AND read_state)) OR ((reconfig_mode_sel(3) AND reconfig_mode_sel(2)) AND reconfig_mode_sel(1))) OR (wire_w99w(0) AND wire_w_lg_write_done91w(0)));
	is_illegal_reg_out <= is_illegal_reg;
	is_pll_address <= '0';
	is_protected_bit <= '0';
	is_rcxpat_chnl_en_ch <= '0';
	is_table_33 <= '0';
	is_table_59 <= '0';
	is_table_61 <= '0';
	is_tier_1 <= '0';
	is_tier_2 <= '0';
	is_tx_local_div_ctrl <= '0';
	local_ch_dec <= wire_aeq_ch_done_mux_result(0);
	logical_pll_sel_num <= (OTHERS => '0');
	mif_family_error <= '0';
	mif_reconfig_done <= '0';
	mif_type_error <= '0';
	offset_cancellation_reset <= '0';
	quad_address <= ( "000" & wire_addr_cntr_q(7 DOWNTO 2));
	quad_address_out <= address_pres_reg(11 DOWNTO 3);
	rate_switch_ctrl_max_limit <= "000000000011";
	rd_pulse <= (((((wire_w_lg_dprio_pulse581w(0) AND wire_w_lg_write_done91w(0)) AND wire_wr_rd_pulse_reg_w_lg_q570w(0)) AND wire_w_lg_write_state596w(0)) OR (wire_w_lg_read_state582w(0) AND wire_w_lg_read_done580w(0))) AND wire_w_lg_is_illegal_reg_d579w(0));
	read_addr_inc <= (read_state AND dprio_pulse);
	read_address <= ( "0" & address_pres_reg(2) & channel_address_out & "1" & wire_read_addr_cntr_q(2) & "000000" & wire_read_addr_cntr_w_lg_w_q_range693w696w & "0" & wire_read_addr_cntr_w_lg_w_q_range699w700w & wire_read_addr_cntr_q(0));
	read_done <= (((read_word_done AND read_addr_inc) OR (is_illegal_reg_out AND read_state)) OR reset_system);
	read_state <= (state_mc_reg(0) AND wire_state_mc_reg_w_lg_q29w(0));
	read_word_64_67_data_valid <= ((wire_w_lg_dprio_pulse716w(0) AND (NOT wire_read_addr_cntr_q(1))) AND (NOT wire_read_addr_cntr_q(0)));
	read_word_68_6B_data_valid <= ((wire_w_lg_dprio_pulse716w(0) AND (NOT wire_read_addr_cntr_q(1))) AND wire_read_addr_cntr_q(0));
	read_word_7c_7f_data_valid <= ((wire_w_lg_dprio_pulse709w(0) AND wire_read_addr_cntr_q(1)) AND (NOT wire_read_addr_cntr_q(0)));
	read_word_7c_7f_inv_data_valid <= ((wire_w_lg_dprio_pulse709w(0) AND wire_read_addr_cntr_q(1)) AND wire_read_addr_cntr_q(0));
	read_word_done <= ((read_word_68_6B_data_valid AND rx_reconfig) OR wire_w_lg_read_word_7c_7f_inv_data_valid703w(0));
	read_word_preemp_1t_data_valid <= ((wire_w_lg_dprio_pulse709w(0) AND (NOT wire_read_addr_cntr_q(1))) AND wire_read_addr_cntr_q(0));
	read_word_vodctrl_data_valid <= ((wire_w_lg_dprio_pulse709w(0) AND (NOT wire_read_addr_cntr_q(1))) AND (NOT wire_read_addr_cntr_q(0)));
	reconfig_datain <= (OTHERS => '0');
	reconfig_reset_all <= '0';
	reconfig_togxb <= ( wire_calibration_busy & wire_dprio_dprioload & wire_dprio_dpriodisable & wire_dprio_dprioin);
	remap_eyemon <= ((wire_w_lg_w_reconfig_mode_sel_range644w645w(0) AND reconfig_mode_sel(2)) AND reconfig_mode_sel(3));
	reset_addr_done <= '0';
	reset_reconf_addr <= '0';
	reset_system <= reset_system_reg;
	rx_eqctrl_out <= rx_eqctrl_reg;
	rx_eqdcgain_out <= rx_equalizer_dcgain_reg;
	rx_reconfig <= '1';
	s0_to_0 <= ((idle_state AND write_all_int) OR read_done);
	s0_to_1 <= ((wire_w_lg_idle_state50w(0) AND wire_w_lg_write_state48w(0)) AND wire_w_lg_write_all_int47w(0));
	s0_to_2 <= (wire_w_lg_idle_state41w(0) AND (wire_w_lg_write_all25w(0) OR (is_bonded_reconfig AND is_bonded_global_clk_div)));
	s1_to_0 <= ((wire_w_lg_idle_state50w(0) AND wire_w_lg_write_state48w(0)) OR write_done);
	s1_to_1 <= (idle_state AND write_all_int);
	s2_to_0 <= (adce_state AND (NOT ((adce_busy_state OR eyemon_busy) OR dfe_busy)));
	sel_max_limit <= ((((wire_w_lg_w_lg_is_analog_control108w109w OR wire_w_lg_w_lg_is_analog_control106w107w) OR wire_w_lg_is_tier_1105w) OR wire_w_lg_is_tx_local_div_ctrl104w) OR wire_w_lg_is_adce_mode_sel103w);
	start <= '0';
	state_mc_reg_in <= ( wire_w_lg_w_lg_s0_to_273w74w & wire_w_lg_w_lg_s0_to_262w63w);
	tier_1_max_limit <= "000000000111";
	transceiver_init <= '0';
	tx_preemp_0t_out <= ( wire_tx_preemp_0t_inv_reg_w_lg_w_q_range1139w1140w & wire_add_sub11_result);
	tx_preemp_0t_out_wire <= tx_preemphasisctrl_pretap_reg;
	tx_preemp_0t_wire <= wire_add_sub1_result;
	tx_preemp_1t_out <= tx_preemphasisctrl_1stposttap_reg;
	tx_preemp_2t_out <= ( wire_tx_preemp_2t_inv_reg_w_lg_w_q_range1149w1150w & wire_add_sub12_result);
	tx_preemp_2t_out_wire <= tx_preemphasisctrl_2ndposttap_reg;
	tx_preemp_2t_wire <= wire_add_sub2_result;
	tx_reconfig <= '1';
	tx_vodctrl_out <= tx_vodctrl_reg;
	wire_w185w <= ( cal_quad_address & cal_channel_address(2 DOWNTO 0));
	w721w <= ( quad_address & channel_address);
	w_eq_0_1004w <= ( "0" & "0" & wire_w_lg_w_w_rx_eqv959w_range1014w1015w & wire_w1024w);
	w_eq_10_1045w <= ( "1" & wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1049w1050w & wire_w1052w & wire_w1055w);
	w_eq_3_1026w <= ( "0" & "1" & wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1022w1023w & wire_w_lg_w_lg_w_w_rx_eqv959w_range1014w1033w1034w);
	w_eq_6_1036w <= ( w_rx_eqv959w(2) & wire_w_lg_w_w_rx_eqv959w_range1014w1019w & wire_w1024w & wire_w_lg_w_lg_w_w_rx_eqv959w_range1011w1018w1043w);
	w_gt_0_964w <= ((w_rx_eqd955w(2) AND w_rx_eqd955w(1)) AND w_rx_eqd955w(0));
	w_gt_0_only988w <= ((wire_w_lg_w_gt_0_964w992w(0) AND wire_w_lg_w_gt_6_976w990w(0)) AND wire_w_lg_w_gt_10_982w989w(0));
	w_gt_10_982w <= ((w_rx_eqa958w(2) AND w_rx_eqa958w(1)) AND w_rx_eqa958w(0));
	w_gt_10_only1002w <= (wire_w_lg_w_lg_w_gt_0_964w996w1000w(0) AND ((w_rx_eqa958w(2) AND w_rx_eqa958w(1)) AND w_rx_eqa958w(0)));
	w_gt_3_970w <= ((w_rx_eqc956w(2) AND w_rx_eqc956w(1)) AND w_rx_eqc956w(0));
	w_gt_3_only995w <= ((wire_w_lg_w_gt_0_964w996w(0) AND wire_w_lg_w_gt_6_976w990w(0)) AND wire_w_lg_w_gt_10_982w989w(0));
	w_gt_6_976w <= ((w_rx_eqb957w(2) AND w_rx_eqb957w(1)) AND w_rx_eqb957w(0));
	w_gt_6_only999w <= (wire_w_lg_w_lg_w_gt_0_964w996w1000w(0) AND wire_w_lg_w_gt_10_982w989w(0));
	w_rx_eqa958w <= wire_dprio_dataout(14 DOWNTO 12);
	w_rx_eqb957w <= wire_dprio_dataout(11 DOWNTO 9);
	w_rx_eqc956w <= wire_dprio_dataout(8 DOWNTO 6);
	w_rx_eqctrl_out954w <= (((wire_w_lg_w_eq_0_1004w1060w OR wire_w_lg_w_eq_3_1026w1059w) OR wire_w_lg_w_eq_6_1036w1058w) OR wire_w_lg_w_eq_10_1045w1057w);
	w_rx_eqd955w <= wire_dprio_dataout(5 DOWNTO 3);
	w_rx_eqdcgain_out1070w <= ( wire_dprio_dataout(10) & wire_dprio_w_lg_w_dataout_range1075w1076w & wire_dprio_w_lg_w_lg_w_lg_w_dataout_range1079w1080w1081w1082w);
	w_rx_eqv959w <= wire_dprio_dataout(2 DOWNTO 0);
	w_tx_vodctrl_out1090w <= ( wire_dprio_w_lg_w_lg_w_dataout_range1091w1095w1096w & wire_dprio_w_lg_w_lg_w_dataout_range1091w1100w1101w & wire_dprio_w_lg_w_lg_w_lg_w_dataout_range1091w1092w1104w1105w);
	w_wire_adce_dprioout_mux2434w <= ( wire_w_lg_w_lg_adce_busy_state132w509w & wire_w_lg_w_lg_adce_busy_state132w497w & wire_w_lg_w_lg_adce_busy_state132w485w & wire_w_lg_w_lg_adce_busy_state132w473w & wire_w_lg_w_lg_adce_busy_state132w461w & wire_w_lg_w_lg_adce_busy_state132w448w);
	w_wire_adce_dprioout_mux433w <= ( wire_w_lg_adce_busy_state506w & wire_w_lg_adce_busy_state494w & wire_w_lg_adce_busy_state482w & wire_w_lg_adce_busy_state470w & wire_w_lg_adce_busy_state458w & wire_w_lg_adce_busy_state444w);
	w_wire_dfe_dprioout_mux431w <= ( wire_w_lg_dfe_busy500w & wire_w_lg_dfe_busy488w & wire_w_lg_dfe_busy476w & wire_w_lg_dfe_busy464w & wire_w_lg_dfe_busy452w & wire_w_lg_dfe_busy436w);
	w_wire_eyemon_dprioout_mux432w <= ( wire_w_lg_eyemon_busy503w & wire_w_lg_eyemon_busy491w & wire_w_lg_eyemon_busy479w & wire_w_lg_eyemon_busy467w & wire_w_lg_eyemon_busy455w & wire_w_lg_eyemon_busy440w);
	wr_pulse <= (((wire_w_lg_write_state619w(0) AND wire_w_lg_write_done91w(0)) AND (wire_wr_rd_pulse_reg_w_lg_q617w(0) OR (wire_w_lg_is_tier_1613w(0) AND (((((wire_w_lg_is_rcxpat_chnl_en_ch607w(0) AND wire_w_lg_is_cruclk_addr0606w(0)) AND wire_w_lg_write_skip605w(0)) AND wire_w_lg_bonded_skip604w(0)) AND wire_w_lg_is_protected_bit603w(0)) AND wire_w_lg_is_global_clk_div_mode602w(0))))) AND wire_w_lg_is_illegal_reg_d579w(0));
	write_addr_inc <= ((write_state AND dprio_pulse) AND write_happened);
	write_address <= ( "0" & address_pres_reg(2) & channel_address_out & "1" & wire_write_addr_cntr_q(2) & "000000" & wire_write_addr_cntr_w_lg_w_q_range928w931w & "0" & wire_write_addr_cntr_w_lg_w_q_range934w935w & wire_write_addr_cntr_q(0));
	write_all_int <= ((wire_w_lg_write_all25w(0) OR (is_bonded_reconfig AND is_bonded_global_clk_div)) AND en_write_trigger);
	write_done <= ((wire_w_lg_w_lg_write_word_done906w907w(0) OR (is_illegal_reg_out AND write_state)) OR reset_system);
	write_happened <= wr_addr_inc_reg;
	write_skip <= '0';
	write_state <= (wire_state_mc_reg_w_lg_q31w(0) AND state_mc_reg(1));
	write_word_64_67_data_valid <= (wire_write_addr_cntr_w_lg_w_q_range928w951w(0) AND (NOT wire_write_addr_cntr_q(0)));
	write_word_68_6B_data_valid <= (wire_write_addr_cntr_w_lg_w_q_range928w951w(0) AND wire_write_addr_cntr_q(0));
	write_word_7c_7f_data_valid <= (((NOT wire_write_addr_cntr_q(2)) AND wire_write_addr_cntr_q(1)) AND (NOT wire_write_addr_cntr_q(0)));
	write_word_7c_7f_inv_data_valid <= (((NOT wire_write_addr_cntr_q(2)) AND wire_write_addr_cntr_q(1)) AND wire_write_addr_cntr_q(0));
	write_word_done <= (dprio_pulse AND ((write_word_68_6B_data_valid AND rx_reconfig) OR wire_w_lg_write_word_7c_7f_inv_data_valid938w(0)));
	write_word_preemp1t_data_valid <= (((NOT wire_write_addr_cntr_q(2)) AND wire_write_addr_cntr_w_lg_w_q_range934w943w(0)) AND wire_write_addr_cntr_q(0));
	write_word_preemp1ta_data_valid <= '0';
	write_word_preemp1tb_data_valid <= '0';
	write_word_vodctrl_data_valid <= (((NOT wire_write_addr_cntr_q(2)) AND wire_write_addr_cntr_w_lg_w_q_range934w943w(0)) AND (NOT wire_write_addr_cntr_q(0)));
	write_word_vodctrla_data_valid <= '0';
	wire_w_adce_quad_addr_s4_range443w(0) <= adce_quad_addr_s4(0);
	wire_w_adce_quad_addr_s4_range457w(0) <= adce_quad_addr_s4(1);
	wire_w_adce_quad_addr_s4_range469w(0) <= adce_quad_addr_s4(2);
	wire_w_adce_quad_addr_s4_range481w(0) <= adce_quad_addr_s4(3);
	wire_w_adce_quad_addr_s4_range493w(0) <= adce_quad_addr_s4(4);
	wire_w_adce_quad_addr_s4_range505w(0) <= adce_quad_addr_s4(5);
	wire_w_cal_quad_address_range515w(0) <= cal_quad_address(0);
	wire_w_cal_quad_address_range524w(0) <= cal_quad_address(1);
	wire_w_cal_quad_address_range532w(0) <= cal_quad_address(2);
	wire_w_cal_quad_address_range540w(0) <= cal_quad_address(3);
	wire_w_cal_quad_address_range548w(0) <= cal_quad_address(4);
	wire_w_cal_quad_address_range556w(0) <= cal_quad_address(5);
	wire_w_channel_address_range153w(0) <= channel_address(0);
	wire_w_channel_address_range143w(0) <= channel_address(1);
	wire_w_dfe_quad_address_range435w(0) <= dfe_quad_address(0);
	wire_w_dfe_quad_address_range451w(0) <= dfe_quad_address(1);
	wire_w_dfe_quad_address_range463w(0) <= dfe_quad_address(2);
	wire_w_dfe_quad_address_range475w(0) <= dfe_quad_address(3);
	wire_w_dfe_quad_address_range487w(0) <= dfe_quad_address(4);
	wire_w_dfe_quad_address_range499w(0) <= dfe_quad_address(5);
	wire_w_eyemon_quad_address_range439w(0) <= eyemon_quad_address(0);
	wire_w_eyemon_quad_address_range454w(0) <= eyemon_quad_address(1);
	wire_w_eyemon_quad_address_range466w(0) <= eyemon_quad_address(2);
	wire_w_eyemon_quad_address_range478w(0) <= eyemon_quad_address(3);
	wire_w_eyemon_quad_address_range490w(0) <= eyemon_quad_address(4);
	wire_w_eyemon_quad_address_range502w(0) <= eyemon_quad_address(5);
	wire_w_logical_pll_sel_num_range150w(0) <= logical_pll_sel_num(0);
	wire_w_logical_pll_sel_num_range139w(0) <= logical_pll_sel_num(1);
	wire_w_quad_address_range447w(0) <= quad_address(0);
	wire_w_quad_address_range460w(0) <= quad_address(1);
	wire_w_quad_address_range472w(0) <= quad_address(2);
	wire_w_quad_address_range484w(0) <= quad_address(3);
	wire_w_quad_address_range496w(0) <= quad_address(4);
	wire_w_quad_address_range508w(0) <= quad_address(5);
	wire_w_reconfig_mode_sel_range644w(0) <= reconfig_mode_sel(0);
	wire_w_reconfig_mode_sel_range85w(0) <= reconfig_mode_sel(1);
	wire_w_rx_eqctrl_range845w(0) <= rx_eqctrl(0);
	wire_w_rx_eqctrl_range838w(0) <= rx_eqctrl(1);
	wire_w_rx_eqctrl_range840w(0) <= rx_eqctrl(2);
	wire_w_rx_eqctrl_range842w(0) <= rx_eqctrl(3);
	wire_w_rx_eqdcgain_range819w(0) <= rx_eqdcgain(0);
	wire_w_rx_eqdcgain_range820w(0) <= rx_eqdcgain(1);
	wire_w_rx_eqdcgain_range816w(0) <= rx_eqdcgain(2);
	wire_w_tx_preemp_0t_range2w(0) <= tx_preemp_0t(4);
	wire_w_tx_preemp_0t_wire_range894w <= tx_preemp_0t_wire(3 DOWNTO 0);
	wire_w_tx_preemp_2t_range4w(0) <= tx_preemp_2t(4);
	wire_w_tx_preemp_2t_wire_range898w <= tx_preemp_2t_wire(3 DOWNTO 0);
	wire_w_tx_vodctrl_range761w(0) <= tx_vodctrl(0);
	wire_w_tx_vodctrl_range758w(0) <= tx_vodctrl(1);
	wire_w_tx_vodctrl_range759w(0) <= tx_vodctrl(2);
	wire_w_w_rx_eqv959w_range1010w(0) <= w_rx_eqv959w(0);
	wire_w_w_rx_eqv959w_range1011w(0) <= w_rx_eqv959w(1);
	wire_w_w_rx_eqv959w_range1014w(0) <= w_rx_eqv959w(2);
	wire_w_w_wire_adce_dprioout_mux2434w_range449w(0) <= w_wire_adce_dprioout_mux2434w(0);
	wire_w_w_wire_adce_dprioout_mux2434w_range462w(0) <= w_wire_adce_dprioout_mux2434w(1);
	wire_w_w_wire_adce_dprioout_mux2434w_range474w(0) <= w_wire_adce_dprioout_mux2434w(2);
	wire_w_w_wire_adce_dprioout_mux2434w_range486w(0) <= w_wire_adce_dprioout_mux2434w(3);
	wire_w_w_wire_adce_dprioout_mux2434w_range498w(0) <= w_wire_adce_dprioout_mux2434w(4);
	wire_w_w_wire_adce_dprioout_mux2434w_range510w(0) <= w_wire_adce_dprioout_mux2434w(5);
	wire_w_w_wire_adce_dprioout_mux433w_range445w(0) <= w_wire_adce_dprioout_mux433w(0);
	wire_w_w_wire_adce_dprioout_mux433w_range459w(0) <= w_wire_adce_dprioout_mux433w(1);
	wire_w_w_wire_adce_dprioout_mux433w_range471w(0) <= w_wire_adce_dprioout_mux433w(2);
	wire_w_w_wire_adce_dprioout_mux433w_range483w(0) <= w_wire_adce_dprioout_mux433w(3);
	wire_w_w_wire_adce_dprioout_mux433w_range495w(0) <= w_wire_adce_dprioout_mux433w(4);
	wire_w_w_wire_adce_dprioout_mux433w_range507w(0) <= w_wire_adce_dprioout_mux433w(5);
	wire_w_w_wire_dfe_dprioout_mux431w_range437w(0) <= w_wire_dfe_dprioout_mux431w(0);
	wire_w_w_wire_dfe_dprioout_mux431w_range453w(0) <= w_wire_dfe_dprioout_mux431w(1);
	wire_w_w_wire_dfe_dprioout_mux431w_range465w(0) <= w_wire_dfe_dprioout_mux431w(2);
	wire_w_w_wire_dfe_dprioout_mux431w_range477w(0) <= w_wire_dfe_dprioout_mux431w(3);
	wire_w_w_wire_dfe_dprioout_mux431w_range489w(0) <= w_wire_dfe_dprioout_mux431w(4);
	wire_w_w_wire_dfe_dprioout_mux431w_range501w(0) <= w_wire_dfe_dprioout_mux431w(5);
	wire_w_w_wire_eyemon_dprioout_mux432w_range441w(0) <= w_wire_eyemon_dprioout_mux432w(0);
	wire_w_w_wire_eyemon_dprioout_mux432w_range456w(0) <= w_wire_eyemon_dprioout_mux432w(1);
	wire_w_w_wire_eyemon_dprioout_mux432w_range468w(0) <= w_wire_eyemon_dprioout_mux432w(2);
	wire_w_w_wire_eyemon_dprioout_mux432w_range480w(0) <= w_wire_eyemon_dprioout_mux432w(3);
	wire_w_w_wire_eyemon_dprioout_mux432w_range492w(0) <= w_wire_eyemon_dprioout_mux432w(4);
	wire_w_w_wire_eyemon_dprioout_mux432w_range504w(0) <= w_wire_eyemon_dprioout_mux432w(5);
	wire_calibration_w_lg_w_lg_busy377w428w(0) <= wire_calibration_w_lg_busy377w(0) AND a2gr_dprio_wren_data;
	loop54 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_w_lg_busy377w391w(i) <= wire_calibration_w_lg_busy377w(0) AND wire_adce_dprio_addr_mux_result(i);
	END GENERATE loop54;
	loop55 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_w_lg_busy377w378w(i) <= wire_calibration_w_lg_busy377w(0) AND wire_adce_dprio_data_mux_result(i);
	END GENERATE loop55;
	loop56 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_busy392w(i) <= wire_calibration_busy AND cal_dprio_address(i);
	END GENERATE loop56;
	loop57 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_busy379w(i) <= wire_calibration_busy AND wire_calibration_dprio_dataout(i);
	END GENERATE loop57;
	wire_calibration_w_lg_busy377w(0) <= NOT wire_calibration_busy;
	wire_calibration_reset <= wire_w_lg_offset_cancellation_reset207w(0);
	wire_w_lg_offset_cancellation_reset207w(0) <= offset_cancellation_reset OR reconfig_reset_all;
	calibration :  alt_cal
	  GENERIC MAP (
		CHANNEL_ADDRESS_WIDTH => 8,
		NUMBER_OF_CHANNELS => 144,
		SIM_MODEL_MODE => "FALSE"
	  )
	  PORT MAP ( 
		busy => wire_calibration_busy,
		clock => reconfig_clk,
		dprio_addr => wire_calibration_dprio_addr,
		dprio_busy => wire_dprio_busy,
		dprio_datain => wire_dprio_dataout,
		dprio_dataout => wire_calibration_dprio_dataout,
		dprio_rden => wire_calibration_dprio_rden,
		dprio_wren => wire_calibration_dprio_wren,
		quad_addr => wire_calibration_quad_addr,
		remap_addr => address_pres_reg,
		reset => wire_calibration_reset,
		retain_addr => wire_calibration_retain_addr,
		start => start,
		testbuses => cal_testbuses,
		transceiver_init => transceiver_init
	  );
	wire_dfe_i_avmm_saddress <= wire_w_lg_ctrl_address365w;
	wire_dfe_i_avmm_sread <= wire_w_lg_ctrl_read366w(0);
	wire_w_lg_ctrl_read366w(0) <= ctrl_read AND wire_w_lg_is_do_eyemon364w(0);
	wire_dfe_i_avmm_swrite <= wire_w_lg_ctrl_write367w(0);
	wire_w_lg_ctrl_write367w(0) <= ctrl_write AND wire_w_lg_is_do_eyemon364w(0);
	wire_dfe_i_avmm_swritedata <= wire_w_lg_ctrl_writedata368w;
	wire_dfe_i_resetn <= wire_w_lg_reconfig_reset_all28w(0);
	dfe :  alt_dfe
	  GENERIC MAP (
		channel_address_width => 8,
		ireg_chaddr_width => 8
	  )
	  PORT MAP ( 
		i_avmm_clk => reconfig_clk,
		i_avmm_saddress => wire_dfe_i_avmm_saddress,
		i_avmm_sread => wire_dfe_i_avmm_sread,
		i_avmm_swrite => wire_dfe_i_avmm_swrite,
		i_avmm_swritedata => wire_dfe_i_avmm_swritedata,
		i_dprio_busy => wire_dprio_busy,
		i_dprio_in => wire_dprio_dataout,
		i_remap_address => address_pres_reg,
		i_resetn => wire_dfe_i_resetn,
		o_avmm_sreaddata => wire_dfe_o_avmm_sreaddata,
		o_avmm_swaitrequest => wire_dfe_o_avmm_swaitrequest,
		o_dprio_addr => wire_dfe_o_dprio_addr,
		o_dprio_data => wire_dfe_o_dprio_data,
		o_dprio_rden => wire_dfe_o_dprio_rden,
		o_dprio_wren => wire_dfe_o_dprio_wren,
		o_quad_address => wire_dfe_o_quad_address,
		o_reconfig_busy => wire_dfe_o_reconfig_busy
	  );
	wire_dprio_w_lg_w_lg_w_dataout_range1091w1092w1104w(0) <= wire_dprio_w_lg_w_dataout_range1091w1092w(0) AND wire_dprio_w_dataout_range1094w(0);
	wire_dprio_w_lg_w_dataout_range1091w1100w(0) <= wire_dprio_w_dataout_range1091w(0) AND wire_dprio_w_lg_w_dataout_range1094w1099w(0);
	wire_dprio_w_lg_w_dataout_range1091w1095w(0) <= wire_dprio_w_dataout_range1091w(0) AND wire_dprio_w_dataout_range1094w(0);
	wire_dprio_w_lg_w_dataout_range884w1093w(0) <= wire_dprio_w_dataout_range884w(0) AND wire_dprio_w_lg_w_dataout_range1091w1092w(0);
	wire_dprio_w_lg_w_dataout_range884w1103w(0) <= wire_dprio_w_dataout_range884w(0) AND wire_dprio_w_dataout_range1091w(0);
	wire_dprio_w_lg_w_dataout_range1075w1076w(0) <= wire_dprio_w_dataout_range1075w(0) AND wire_dprio_w_lg_w_dataout_range1071w1074w(0);
	wire_dprio_w_lg_busy567w(0) <= NOT wire_dprio_busy;
	wire_dprio_w_lg_w_dataout_range1071w1074w(0) <= NOT wire_dprio_w_dataout_range1071w(0);
	wire_dprio_w_lg_w_dataout_range1094w1099w(0) <= NOT wire_dprio_w_dataout_range1094w(0);
	wire_dprio_w_lg_w_dataout_range1091w1092w(0) <= NOT wire_dprio_w_dataout_range1091w(0);
	wire_dprio_w_lg_w_lg_w_lg_w_dataout_range1091w1092w1104w1105w(0) <= wire_dprio_w_lg_w_lg_w_dataout_range1091w1092w1104w(0) OR wire_dprio_w_lg_w_dataout_range884w1103w(0);
	wire_dprio_w_lg_w_lg_w_dataout_range1091w1100w1101w(0) <= wire_dprio_w_lg_w_dataout_range1091w1100w(0) OR wire_dprio_w_lg_w_dataout_range884w1093w(0);
	wire_dprio_w_lg_w_lg_w_dataout_range1091w1095w1096w(0) <= wire_dprio_w_lg_w_dataout_range1091w1095w(0) OR wire_dprio_w_lg_w_dataout_range884w1093w(0);
	wire_dprio_w_lg_w_lg_w_lg_w_dataout_range1079w1080w1081w1082w(0) <= wire_dprio_w_lg_w_lg_w_dataout_range1079w1080w1081w(0) XOR wire_dprio_w_dataout_range1071w(0);
	wire_dprio_w_lg_w_lg_w_dataout_range1079w1080w1081w(0) <= wire_dprio_w_lg_w_dataout_range1079w1080w(0) XOR wire_dprio_w_dataout_range1078w(0);
	wire_dprio_w_lg_w_dataout_range1079w1080w(0) <= wire_dprio_w_dataout_range1079w(0) XOR wire_dprio_w_dataout_range1075w(0);
	wire_dprio_address <= wire_calibration_w_lg_w_lg_busy392w393w;
	loop58 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_w_lg_busy392w393w(i) <= wire_calibration_w_lg_busy392w(i) OR wire_calibration_w_lg_w_lg_busy377w391w(i);
	END GENERATE loop58;
	wire_dprio_datain <= wire_calibration_w_lg_w_lg_busy379w380w;
	loop59 : FOR i IN 0 TO 15 GENERATE 
		wire_calibration_w_lg_w_lg_busy379w380w(i) <= wire_calibration_w_lg_busy379w(i) OR wire_calibration_w_lg_w_lg_busy377w378w(i);
	END GENERATE loop59;
	wire_dprio_rden <= wire_calibration_w_lg_w_lg_busy413w414w(0);
	wire_calibration_w_lg_w_lg_busy413w414w(0) <= (wire_calibration_busy AND wire_calibration_dprio_rden) OR (wire_calibration_w_lg_busy377w(0) AND wire_adce_dprio_enas_mux_result(0));
	wire_dprio_wren <= wire_calibration_w_lg_w_lg_busy417w418w(0);
	wire_calibration_w_lg_w_lg_busy417w418w(0) <= (wire_calibration_busy AND wire_calibration_dprio_wren) OR (wire_calibration_w_lg_busy377w(0) AND wire_adce_dprio_enas_mux_result(1));
	wire_dprio_wren_data <= wire_calibration_w_lg_w_lg_busy429w430w(0);
	wire_calibration_w_lg_w_lg_busy429w430w(0) <= (wire_calibration_busy AND wire_calibration_retain_addr) OR wire_calibration_w_lg_w_lg_busy377w428w(0);
	wire_dprio_w_dataout_range1071w(0) <= wire_dprio_dataout(10);
	wire_dprio_w_dataout_range1094w(0) <= wire_dprio_dataout(13);
	wire_dprio_w_dataout_range1091w(0) <= wire_dprio_dataout(14);
	wire_dprio_w_dataout_range797w <= wire_dprio_dataout(15 DOWNTO 11);
	wire_dprio_w_dataout_range884w(0) <= wire_dprio_dataout(15);
	wire_dprio_w_dataout_range1117w <= wire_dprio_dataout(3 DOWNTO 0);
	wire_dprio_w_dataout_range1136w(0) <= wire_dprio_dataout(4);
	wire_dprio_w_dataout_range1129w <= wire_dprio_dataout(7 DOWNTO 4);
	wire_dprio_w_dataout_range1079w(0) <= wire_dprio_dataout(7);
	wire_dprio_w_dataout_range1075w(0) <= wire_dprio_dataout(8);
	wire_dprio_w_dataout_range1078w(0) <= wire_dprio_dataout(9);
	wire_dprio_w_dataout_range1146w(0) <= wire_dprio_dataout(3);
	dprio :  reconfig_side_alt_dprio_2vj
	  PORT MAP ( 
		address => wire_dprio_address,
		busy => wire_dprio_busy,
		datain => wire_dprio_datain,
		dataout => wire_dprio_dataout,
		dpclk => reconfig_clk,
		dpriodisable => wire_dprio_dpriodisable,
		dprioin => wire_dprio_dprioin,
		dprioload => wire_dprio_dprioload,
		dprioout => wire_dprioout_mux_result(0),
		quad_address => quad_address_out,
		rden => wire_dprio_rden,
		reset => reconfig_reset_all,
		wren => wire_dprio_wren,
		wren_data => wire_dprio_wren_data
	  );
	wire_eyemonitor_i_avmm_saddress <= wire_w_lg_ctrl_address357w;
	wire_eyemonitor_i_avmm_sread <= wire_w_lg_ctrl_read358w(0);
	wire_w_lg_ctrl_read358w(0) <= ctrl_read AND wire_w_lg_is_do_dfe356w(0);
	wire_eyemonitor_i_avmm_swrite <= wire_w_lg_ctrl_write359w(0);
	wire_w_lg_ctrl_write359w(0) <= ctrl_write AND wire_w_lg_is_do_dfe356w(0);
	wire_eyemonitor_i_avmm_swritedata <= wire_w_lg_ctrl_writedata360w;
	wire_eyemonitor_i_resetn <= wire_w_lg_reconfig_reset_all28w(0);
	eyemonitor :  alt_eyemon
	  GENERIC MAP (
		channel_address_width => 8,
		ireg_chaddr_width => 8
	  )
	  PORT MAP ( 
		i_avmm_clk => reconfig_clk,
		i_avmm_saddress => wire_eyemonitor_i_avmm_saddress,
		i_avmm_sread => wire_eyemonitor_i_avmm_sread,
		i_avmm_swrite => wire_eyemonitor_i_avmm_swrite,
		i_avmm_swritedata => wire_eyemonitor_i_avmm_swritedata,
		i_dprio_busy => wire_dprio_busy,
		i_dprio_in => wire_dprio_dataout,
		i_remap_address => address_pres_reg,
		i_remap_phase => remap_eyemon,
		i_resetn => wire_eyemonitor_i_resetn,
		o_avmm_sreaddata => wire_eyemonitor_o_avmm_sreaddata,
		o_avmm_swaitrequest => wire_eyemonitor_o_avmm_swaitrequest,
		o_dprio_addr => wire_eyemonitor_o_dprio_addr,
		o_dprio_data => wire_eyemonitor_o_dprio_data,
		o_dprio_rden => wire_eyemonitor_o_dprio_rden,
		o_dprio_wren => wire_eyemonitor_o_dprio_wren,
		o_quad_address => wire_eyemonitor_o_quad_address,
		o_reconfig_busy => wire_eyemonitor_o_reconfig_busy
	  );
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN address_pres_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN address_pres_reg <= wire_w_lg_w_lg_cal_busy186w187w;
		END IF;
	END PROCESS;
	wire_address_pres_reg_w_lg_w_lg_w_q_range191w192w193w(0) <= wire_address_pres_reg_w_lg_w_q_range191w192w(0) AND wire_address_pres_reg_w_q_range189w(0);
	loop60 : FOR i IN 0 TO 1 GENERATE 
		wire_address_pres_reg_w_lg_w_q_range195w196w(i) <= wire_address_pres_reg_w_q_range195w(i) AND wire_address_pres_reg_w_lg_w_lg_w_lg_w_q_range191w192w193w194w(0);
	END GENERATE loop60;
	wire_address_pres_reg_w_lg_w_q_range191w192w(0) <= wire_address_pres_reg_w_q_range191w(0) AND wire_address_pres_reg_w_q_range190w(0);
	wire_address_pres_reg_w_lg_w_lg_w_lg_w_q_range191w192w193w194w(0) <= NOT wire_address_pres_reg_w_lg_w_lg_w_q_range191w192w193w(0);
	wire_address_pres_reg_w_q_range189w(0) <= address_pres_reg(0);
	wire_address_pres_reg_w_q_range195w <= address_pres_reg(1 DOWNTO 0);
	wire_address_pres_reg_w_q_range190w(0) <= address_pres_reg(1);
	wire_address_pres_reg_w_q_range191w(0) <= address_pres_reg(2);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN data_valid_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_data_valid_reg_ena = '1') THEN data_valid_reg <= (NOT (is_illegal_reg_out OR reset_system));
			END IF;
		END IF;
	END PROCESS;
	wire_data_valid_reg_ena <= (read_state OR write_state);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN dprio_pulse_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_dprio_pulse_reg_ena = '1') THEN dprio_pulse_reg <= wire_dprio_busy;
			END IF;
		END IF;
	END PROCESS;
	wire_dprio_pulse_reg_ena <= (read_state OR write_state);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN error_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN error_reg <= ((is_illegal_reg OR reset_system) OR adce_error_wire);
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN is_illegal_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN is_illegal_reg <= (((wire_w_lg_is_illegal_reg_d124w(0) AND wire_w_lg_is_illegal_reg_out122w(0)) OR wire_w_lg_is_illegal_reg_out121w(0)) OR reset_system);
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reconf_mode_sel_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN reconf_mode_sel_reg <= reconfig_mode_sel;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN reset_system_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
				IF (wire_reset_system_reg_sclr = '1') THEN reset_system_reg <= '0';
				ELSE reset_system_reg <= (wire_max_oper_limit_w_lg_aeb118w(0) AND wire_w_lg_is_adce116w(0));
				END IF;
		END IF;
	END PROCESS;
	wire_reset_system_reg_sclr <= ((mif_reconfig_done OR reset_addr_done) OR is_illegal_reg_out);
	PROCESS (reconfig_clk)
	BEGIN
		IF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_rx_eqctrl_reg_ena(0) = '1') THEN rx_eqctrl_reg(0) <= wire_rx_eqctrl_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk)
	BEGIN
		IF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_rx_eqctrl_reg_ena(1) = '1') THEN rx_eqctrl_reg(1) <= wire_rx_eqctrl_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk)
	BEGIN
		IF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_rx_eqctrl_reg_ena(2) = '1') THEN rx_eqctrl_reg(2) <= wire_rx_eqctrl_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk)
	BEGIN
		IF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_rx_eqctrl_reg_ena(3) = '1') THEN rx_eqctrl_reg(3) <= wire_rx_eqctrl_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	wire_rx_eqctrl_reg_d <= wire_w_lg_w_lg_read_state1068w1069w;
	loop61 : FOR i IN 0 TO 3 GENERATE
		wire_rx_eqctrl_reg_ena(i) <= wire_w_lg_w_lg_read_word_68_6B_data_valid1065w1066w(0);
	END GENERATE loop61;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN rx_equalizer_dcgain_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_rx_equalizer_dcgain_reg_ena(0) = '1') THEN rx_equalizer_dcgain_reg(0) <= wire_rx_equalizer_dcgain_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN rx_equalizer_dcgain_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_rx_equalizer_dcgain_reg_ena(1) = '1') THEN rx_equalizer_dcgain_reg(1) <= wire_rx_equalizer_dcgain_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN rx_equalizer_dcgain_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_rx_equalizer_dcgain_reg_ena(2) = '1') THEN rx_equalizer_dcgain_reg(2) <= wire_rx_equalizer_dcgain_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	wire_rx_equalizer_dcgain_reg_d <= wire_w_lg_w_lg_read_state1088w1089w;
	loop62 : FOR i IN 0 TO 2 GENERATE
		wire_rx_equalizer_dcgain_reg_ena(i) <= wire_w_lg_w_lg_read_word_64_67_data_valid1085w1086w(0);
	END GENERATE loop62;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN state_mc_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN state_mc_reg <= state_mc_reg_in;
		END IF;
	END PROCESS;
	wire_state_mc_reg_w_lg_q31w(0) <= NOT state_mc_reg(0);
	wire_state_mc_reg_w_lg_q29w(0) <= NOT state_mc_reg(1);
	wire_state_mc_reg_w_q_range55w(0) <= state_mc_reg(0);
	wire_state_mc_reg_w_q_range67w(0) <= state_mc_reg(1);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemp_0t_inv_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemp_0t_inv_reg_ena = "1") THEN tx_preemp_0t_inv_reg(0) <= (wire_w_lg_read_state1137w(0) OR wire_w_lg_write_state1135w(0));
			END IF;
		END IF;
	END PROCESS;
	wire_tx_preemp_0t_inv_reg_ena(0) <= ((read_word_7c_7f_inv_data_valid AND read_state) OR (write_state AND write_word_7c_7f_inv_data_valid));
	wire_tx_preemp_0t_inv_reg_w_lg_w_q_range1139w1140w(0) <= NOT wire_tx_preemp_0t_inv_reg_w_q_range1139w(0);
	wire_tx_preemp_0t_inv_reg_w_q_range1139w(0) <= tx_preemp_0t_inv_reg(0);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemp_2t_inv_reg <= (OTHERS => '0');
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemp_2t_inv_reg_ena = "1") THEN tx_preemp_2t_inv_reg(0) <= (wire_w_lg_read_state1147w(0) OR wire_w_lg_write_state1145w(0));
			END IF;
		END IF;
	END PROCESS;
	wire_tx_preemp_2t_inv_reg_ena(0) <= ((read_word_7c_7f_inv_data_valid AND read_state) OR (write_state AND write_word_7c_7f_inv_data_valid));
	wire_tx_preemp_2t_inv_reg_w_lg_w_q_range1149w1150w(0) <= NOT wire_tx_preemp_2t_inv_reg_w_q_range1149w(0);
	wire_tx_preemp_2t_inv_reg_w_q_range1149w(0) <= tx_preemp_2t_inv_reg(0);
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_1stposttap_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_1stposttap_reg_ena(0) = '1') THEN tx_preemphasisctrl_1stposttap_reg(0) <= wire_tx_preemphasisctrl_1stposttap_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_1stposttap_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_1stposttap_reg_ena(1) = '1') THEN tx_preemphasisctrl_1stposttap_reg(1) <= wire_tx_preemphasisctrl_1stposttap_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_1stposttap_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_1stposttap_reg_ena(2) = '1') THEN tx_preemphasisctrl_1stposttap_reg(2) <= wire_tx_preemphasisctrl_1stposttap_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_1stposttap_reg(3) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_1stposttap_reg_ena(3) = '1') THEN tx_preemphasisctrl_1stposttap_reg(3) <= wire_tx_preemphasisctrl_1stposttap_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_1stposttap_reg(4) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_1stposttap_reg_ena(4) = '1') THEN tx_preemphasisctrl_1stposttap_reg(4) <= wire_tx_preemphasisctrl_1stposttap_reg_d(4);
			END IF;
		END IF;
	END PROCESS;
	wire_tx_preemphasisctrl_1stposttap_reg_d <= wire_w_lg_w_lg_read_state1124w1125w;
	loop63 : FOR i IN 0 TO 4 GENERATE
		wire_tx_preemphasisctrl_1stposttap_reg_ena(i) <= wire_w_lg_w_lg_read_word_preemp_1t_data_valid1121w1122w(0);
	END GENERATE loop63;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_2ndposttap_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_2ndposttap_reg_ena(0) = '1') THEN tx_preemphasisctrl_2ndposttap_reg(0) <= wire_tx_preemphasisctrl_2ndposttap_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_2ndposttap_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_2ndposttap_reg_ena(1) = '1') THEN tx_preemphasisctrl_2ndposttap_reg(1) <= wire_tx_preemphasisctrl_2ndposttap_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_2ndposttap_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_2ndposttap_reg_ena(2) = '1') THEN tx_preemphasisctrl_2ndposttap_reg(2) <= wire_tx_preemphasisctrl_2ndposttap_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_2ndposttap_reg(3) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_2ndposttap_reg_ena(3) = '1') THEN tx_preemphasisctrl_2ndposttap_reg(3) <= wire_tx_preemphasisctrl_2ndposttap_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	wire_tx_preemphasisctrl_2ndposttap_reg_d <= wire_w_lg_w_lg_read_state1130w1131w;
	loop64 : FOR i IN 0 TO 3 GENERATE
		wire_tx_preemphasisctrl_2ndposttap_reg_ena(i) <= wire_w_lg_w_lg_read_word_7c_7f_data_valid1126w1127w(0);
	END GENERATE loop64;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_pretap_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_pretap_reg_ena(0) = '1') THEN tx_preemphasisctrl_pretap_reg(0) <= wire_tx_preemphasisctrl_pretap_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_pretap_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_pretap_reg_ena(1) = '1') THEN tx_preemphasisctrl_pretap_reg(1) <= wire_tx_preemphasisctrl_pretap_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_pretap_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_pretap_reg_ena(2) = '1') THEN tx_preemphasisctrl_pretap_reg(2) <= wire_tx_preemphasisctrl_pretap_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_preemphasisctrl_pretap_reg(3) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_preemphasisctrl_pretap_reg_ena(3) = '1') THEN tx_preemphasisctrl_pretap_reg(3) <= wire_tx_preemphasisctrl_pretap_reg_d(3);
			END IF;
		END IF;
	END PROCESS;
	wire_tx_preemphasisctrl_pretap_reg_d <= wire_w_lg_w_lg_read_state1118w1119w;
	loop65 : FOR i IN 0 TO 3 GENERATE
		wire_tx_preemphasisctrl_pretap_reg_ena(i) <= wire_w_lg_w_lg_read_state1114w1115w(0);
	END GENERATE loop65;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_vodctrl_reg(0) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_vodctrl_reg_ena(0) = '1') THEN tx_vodctrl_reg(0) <= wire_tx_vodctrl_reg_d(0);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_vodctrl_reg(1) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_vodctrl_reg_ena(1) = '1') THEN tx_vodctrl_reg(1) <= wire_tx_vodctrl_reg_d(1);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN tx_vodctrl_reg(2) <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_tx_vodctrl_reg_ena(2) = '1') THEN tx_vodctrl_reg(2) <= wire_tx_vodctrl_reg_d(2);
			END IF;
		END IF;
	END PROCESS;
	wire_tx_vodctrl_reg_d <= wire_w_lg_w_lg_read_state1111w1112w;
	loop66 : FOR i IN 0 TO 2 GENERATE
		wire_tx_vodctrl_reg_ena(i) <= wire_w_lg_w_lg_read_word_vodctrl_data_valid1108w1109w(0);
	END GENERATE loop66;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN wr_addr_inc_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN wr_addr_inc_reg <= (wr_pulse OR ((wire_w_lg_wr_pulse199w(0) AND wire_w_lg_rd_pulse198w(0)) AND wr_addr_inc_reg));
		END IF;
	END PROCESS;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN wr_rd_pulse_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_wr_rd_pulse_reg_ena = '1') THEN 
				IF (wire_wr_rd_pulse_reg_sclr = '1') THEN wr_rd_pulse_reg <= '0';
				ELSE wr_rd_pulse_reg <= wire_wr_rd_pulse_reg_w_lg_q570w(0);
				END IF;
			END IF;
		END IF;
	END PROCESS;
	wire_wr_rd_pulse_reg_ena <= (dprio_pulse AND wire_w_lg_read_state571w(0));
	wire_wr_rd_pulse_reg_sclr <= (((wire_w_lg_reset_system575w(0) OR (is_diff_mif AND write_done)) OR reset_addr_done) OR is_illegal_reg_out);
	wire_wr_rd_pulse_reg_w_lg_q617w(0) <= wr_rd_pulse_reg AND wire_w_lg_w_lg_is_tier_1590w616w(0);
	wire_wr_rd_pulse_reg_w_lg_q570w(0) <= NOT wr_rd_pulse_reg;
	PROCESS (reconfig_clk, reconfig_reset_all)
	BEGIN
		IF (reconfig_reset_all = '1') THEN wren_data_reg <= '0';
		ELSIF (reconfig_clk = '1' AND reconfig_clk'event) THEN 
			IF (wire_wren_data_reg_ena = '1') THEN wren_data_reg <= (wire_wren_data_reg_w_lg_w_lg_q724w725w(0) OR wire_wren_data_reg_w_lg_q723w(0));
			END IF;
		END IF;
	END PROCESS;
	wire_wren_data_reg_ena <= (is_tier_1 AND (wire_w_lg_is_diff_mif564w(0) OR (is_diff_mif AND diff_mif_wr_rd_busy)));
	wire_wren_data_reg_w_lg_w_lg_q724w725w(0) <= wire_wren_data_reg_w_lg_q724w(0) AND rd_pulse;
	wire_wren_data_reg_w_lg_q723w(0) <= wren_data_reg AND wire_w_lg_write_done91w(0);
	wire_wren_data_reg_w_lg_q724w(0) <= NOT wren_data_reg;
	wire_wren_data_reg_w_lg_q728w(0) <= wren_data_reg OR is_analog_control;
	wire_add_sub1_dataa <= (OTHERS => '0');
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		add_sub => tx_preemp_0t(4),
		dataa => wire_add_sub1_dataa,
		datab => tx_preemp_0t(3 DOWNTO 0),
		result => wire_add_sub1_result
	  );
	wire_add_sub11_add_sub <= wire_tx_preemp_0t_inv_reg_w_lg_w_q_range1139w1140w(0);
	wire_add_sub11_dataa <= (OTHERS => '0');
	add_sub11 :  lpm_add_sub
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		add_sub => wire_add_sub11_add_sub,
		dataa => wire_add_sub11_dataa,
		datab => tx_preemp_0t_out_wire(3 DOWNTO 0),
		result => wire_add_sub11_result
	  );
	wire_add_sub12_add_sub <= wire_tx_preemp_2t_inv_reg_w_lg_w_q_range1149w1150w(0);
	wire_add_sub12_dataa <= (OTHERS => '0');
	add_sub12 :  lpm_add_sub
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		add_sub => wire_add_sub12_add_sub,
		dataa => wire_add_sub12_dataa,
		datab => tx_preemp_2t_out_wire(3 DOWNTO 0),
		result => wire_add_sub12_result
	  );
	wire_add_sub2_dataa <= (OTHERS => '0');
	add_sub2 :  lpm_add_sub
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		add_sub => tx_preemp_2t(4),
		dataa => wire_add_sub2_dataa,
		datab => tx_preemp_2t(3 DOWNTO 0),
		result => wire_add_sub2_result
	  );
	wire_cmpr10_datab <= (OTHERS => '0');
	cmpr10 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		agb => wire_cmpr10_agb,
		dataa => rx_eqctrl(3 DOWNTO 0),
		datab => wire_cmpr10_datab
	  );
	wire_cmpr7_datab <= "1010";
	cmpr7 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		agb => wire_cmpr7_agb,
		dataa => rx_eqctrl(3 DOWNTO 0),
		datab => wire_cmpr7_datab
	  );
	wire_cmpr8_datab <= "0110";
	cmpr8 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		agb => wire_cmpr8_agb,
		dataa => rx_eqctrl(3 DOWNTO 0),
		datab => wire_cmpr8_datab
	  );
	wire_cmpr9_datab <= "0011";
	cmpr9 :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		agb => wire_cmpr9_agb,
		dataa => rx_eqctrl(3 DOWNTO 0),
		datab => wire_cmpr9_datab
	  );
	wire_max_oper_limit_w_lg_aeb118w(0) <= wire_max_oper_limit_aeb AND wire_w_lg_idle_state117w(0);
	max_oper_limit :  lpm_compare
	  GENERIC MAP (
		LPM_WIDTH => 12
	  )
	  PORT MAP ( 
		aeb => wire_max_oper_limit_aeb,
		dataa => wire_oper_count_q,
		datab => sel_max_limit
	  );
	wire_addr_cntr_sclr <= wire_w_lg_write_done623w(0);
	wire_w_lg_write_done623w(0) <= write_done OR reconfig_reset_all;
	wire_addr_cntr_sload <= wire_w_lg_idle_state625w(0);
	wire_w_lg_idle_state625w(0) <= idle_state AND (write_all OR read);
	addr_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_modulus => 144,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 8
	  )
	  PORT MAP ( 
		clock => reconfig_clk,
		cnt_en => wire_gnd,
		data => logical_channel_address,
		q => wire_addr_cntr_q,
		sclr => wire_addr_cntr_sclr,
		sload => wire_addr_cntr_sload
	  );
	wire_oper_count_sclr <= wire_w_lg_idle_state102w(0);
	wire_w_lg_idle_state102w(0) <= idle_state OR reconfig_reset_all;
	oper_count :  lpm_counter
	  GENERIC MAP (
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 12
	  )
	  PORT MAP ( 
		clock => reconfig_clk,
		cnt_en => dprio_pulse,
		q => wire_oper_count_q,
		sclr => wire_oper_count_sclr
	  );
	wire_read_addr_cntr_w_lg_w_q_range695w698w(0) <= wire_read_addr_cntr_w_q_range695w(0) AND wire_read_addr_cntr_w_q_range693w(0);
	wire_read_addr_cntr_w_lg_w_q_range693w696w(0) <= wire_read_addr_cntr_w_q_range693w(0) AND wire_read_addr_cntr_w_q_range695w(0);
	wire_read_addr_cntr_w_lg_w_q_range693w708w(0) <= NOT wire_read_addr_cntr_w_q_range693w(0);
	wire_read_addr_cntr_w_lg_w_q_range699w700w(0) <= wire_read_addr_cntr_w_q_range699w(0) OR wire_read_addr_cntr_w_lg_w_q_range695w698w(0);
	wire_read_addr_cntr_cnt_en <= wire_w_lg_read_addr_inc674w(0);
	wire_w_lg_read_addr_inc674w(0) <= read_addr_inc AND is_analog_control;
	wire_read_addr_cntr_data <= ( wire_w_lg_tx_reconfig93w & "0" & "0");
	wire_read_addr_cntr_sclr <= wire_w_lg_w_lg_read_done675w676w(0);
	wire_w_lg_w_lg_read_done675w676w(0) <= (read_done OR reset_system) OR reconfig_reset_all;
	wire_read_addr_cntr_sload <= wire_w_lg_w_lg_idle_state683w684w(0);
	wire_w_lg_w_lg_idle_state683w684w(0) <= (idle_state AND read) AND wire_w_lg_tx_reconfig93w(0);
	wire_read_addr_cntr_w_q_range695w(0) <= wire_read_addr_cntr_q(0);
	wire_read_addr_cntr_w_q_range699w(0) <= wire_read_addr_cntr_q(1);
	wire_read_addr_cntr_w_q_range693w(0) <= wire_read_addr_cntr_q(2);
	read_addr_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_modulus => 6,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 3
	  )
	  PORT MAP ( 
		clock => reconfig_clk,
		cnt_en => wire_read_addr_cntr_cnt_en,
		data => wire_read_addr_cntr_data,
		q => wire_read_addr_cntr_q,
		sclr => wire_read_addr_cntr_sclr,
		sload => wire_read_addr_cntr_sload
	  );
	wire_write_addr_cntr_w_lg_w_q_range930w933w(0) <= wire_write_addr_cntr_w_q_range930w(0) AND wire_write_addr_cntr_w_q_range928w(0);
	wire_write_addr_cntr_w_lg_w_q_range928w951w(0) <= wire_write_addr_cntr_w_q_range928w(0) AND wire_write_addr_cntr_w_lg_w_q_range934w943w(0);
	wire_write_addr_cntr_w_lg_w_q_range928w931w(0) <= wire_write_addr_cntr_w_q_range928w(0) AND wire_write_addr_cntr_w_q_range930w(0);
	wire_write_addr_cntr_w_lg_w_q_range934w943w(0) <= NOT wire_write_addr_cntr_w_q_range934w(0);
	wire_write_addr_cntr_w_lg_w_q_range934w935w(0) <= wire_write_addr_cntr_w_q_range934w(0) OR wire_write_addr_cntr_w_lg_w_q_range930w933w(0);
	wire_write_addr_cntr_data <= ( wire_w_lg_tx_reconfig93w & "0" & "0");
	wire_write_addr_cntr_sclr <= wire_w_lg_w_lg_write_done910w911w(0);
	wire_w_lg_w_lg_write_done910w911w(0) <= (write_done OR reset_system) OR reconfig_reset_all;
	wire_write_addr_cntr_sload <= wire_w_lg_w_lg_idle_state918w919w(0);
	wire_w_lg_w_lg_idle_state918w919w(0) <= (idle_state AND write_all) AND wire_w_lg_tx_reconfig93w(0);
	wire_write_addr_cntr_w_q_range930w(0) <= wire_write_addr_cntr_q(0);
	wire_write_addr_cntr_w_q_range934w(0) <= wire_write_addr_cntr_q(1);
	wire_write_addr_cntr_w_q_range928w(0) <= wire_write_addr_cntr_q(2);
	write_addr_cntr :  lpm_counter
	  GENERIC MAP (
		lpm_modulus => 6,
		lpm_port_updown => "PORT_UNUSED",
		lpm_width => 3
	  )
	  PORT MAP ( 
		clock => reconfig_clk,
		cnt_en => write_addr_inc,
		data => wire_write_addr_cntr_data,
		q => wire_write_addr_cntr_q,
		sclr => wire_write_addr_cntr_sclr,
		sload => wire_write_addr_cntr_sload
	  );
	chl_addr_decode :  lpm_decode
	  GENERIC MAP (
		LPM_DECODES => 144,
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		data => wire_addr_cntr_q,
		eq => wire_chl_addr_decode_eq
	  );
	reconf_mode_dec :  lpm_decode
	  GENERIC MAP (
		LPM_DECODES => 16,
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		data => reconf_mode_sel_reg,
		eq => wire_reconf_mode_dec_eq
	  );
	wire_adce_dprio_addr_mux_data <= ( ( eyemon_dprio_addr(15) & address_pres_reg(2) & channel_address_out & eyemon_dprio_addr(11 DOWNTO 0)) & ( dfe_dprio_addr(15 DOWNTO 14) & channel_address_out & dfe_dprio_addr(11 DOWNTO 0)) & ( adce_dprio_addr_s4(15 DOWNTO 14) & channel_address_out & adce_dprio_addr_s4(11 DOWNTO 0)) & a2gr_dprio_addr);
	wire_adce_dprio_addr_mux_sel <= ( wire_w_lg_w_lg_adce_busy_state132w133w & wire_w_lg_adce_busy_state128w);
	adce_dprio_addr_mux :  reconfig_side_mux_t7a
	  PORT MAP ( 
		data => wire_adce_dprio_addr_mux_data,
		result => wire_adce_dprio_addr_mux_result,
		sel => wire_adce_dprio_addr_mux_sel
	  );
	wire_adce_dprio_data_mux_data <= ( eyemon_dprio_data & dfe_dprio_data & adce_dprio_data & a2gr_dprio_data);
	wire_adce_dprio_data_mux_sel <= ( wire_w_lg_w_lg_adce_busy_state132w133w & wire_w_lg_adce_busy_state128w);
	adce_dprio_data_mux :  reconfig_side_mux_t7a
	  PORT MAP ( 
		data => wire_adce_dprio_data_mux_data,
		result => wire_adce_dprio_data_mux_result,
		sel => wire_adce_dprio_data_mux_sel
	  );
	wire_adce_dprio_enas_mux_data <= ( eyemon_dprio_wren & eyemon_dprio_rden & dfe_dprio_wren & dfe_dprio_rden & adce_dprio_wren & adce_dprio_rden & a2gr_dprio_wren & a2gr_dprio_rden);
	wire_adce_dprio_enas_mux_sel <= ( wire_w_lg_w_lg_adce_busy_state132w133w & wire_w_lg_adce_busy_state128w);
	adce_dprio_enas_mux :  reconfig_side_mux_86a
	  PORT MAP ( 
		data => wire_adce_dprio_enas_mux_data,
		result => wire_adce_dprio_enas_mux_result,
		sel => wire_adce_dprio_enas_mux_sel
	  );
	wire_address_pres_reg_mux_data <= ( ( eyemon_pres_reg(11 DOWNTO 0)) & ( dfe_pres_reg(11 DOWNTO 0)) & ( adce_pres_reg(11 DOWNTO 0)) & ( quad_address & wire_w_lg_w_lg_is_pll_address135w136w & wire_w_lg_w146w147w & wire_w_lg_w_lg_w156w157w158w));
	wire_address_pres_reg_mux_sel <= ( wire_w_lg_w_lg_adce_busy_state132w133w & wire_w_lg_adce_busy_state128w);
	address_pres_reg_mux :  reconfig_side_mux_p7a
	  PORT MAP ( 
		data => wire_address_pres_reg_mux_data,
		result => wire_address_pres_reg_mux_result,
		sel => wire_address_pres_reg_mux_sel
	  );
	aeq_ch_done_mux :  reconfig_side_mux_i9a
	  PORT MAP ( 
		data => aeq_ch_done,
		result => wire_aeq_ch_done_mux_result,
		sel => w721w(7 DOWNTO 0)
	  );
	wire_dprioout_mux_sel <= ( wire_w_lg_w_lg_cal_busy557w558w & wire_w_lg_w_lg_cal_busy549w550w & wire_w_lg_w_lg_cal_busy541w542w & wire_w_lg_w_lg_cal_busy533w534w & wire_w_lg_w_lg_cal_busy525w526w & wire_w_lg_w_lg_cal_busy516w517w);
	dprioout_mux :  reconfig_side_mux_08a
	  PORT MAP ( 
		data => cal_dprioout_wire,
		result => wire_dprioout_mux_result,
		sel => wire_dprioout_mux_sel
	  );

 END RTL; --reconfig_side_alt2gxb_reconfig_4og2
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY reconfig_side IS
	PORT
	(
		ctrl_address		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		ctrl_read		: IN STD_LOGIC ;
		ctrl_write		: IN STD_LOGIC ;
		ctrl_writedata		: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		logical_channel_address		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		read		: IN STD_LOGIC ;
		reconfig_clk		: IN STD_LOGIC ;
		reconfig_fromgxb		: IN STD_LOGIC_VECTOR (611 DOWNTO 0);
		reconfig_mode_sel		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		rx_eqctrl		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		rx_eqdcgain		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		tx_preemp_0t		: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		tx_preemp_1t		: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		tx_preemp_2t		: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
		tx_vodctrl		: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
		write_all		: IN STD_LOGIC ;
		busy		: OUT STD_LOGIC ;
		ctrl_readdata		: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		ctrl_waitrequest		: OUT STD_LOGIC ;
		data_valid		: OUT STD_LOGIC ;
		error		: OUT STD_LOGIC ;
		reconfig_togxb		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		rx_eqctrl_out		: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		rx_eqdcgain_out		: OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		tx_preemp_0t_out		: OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
		tx_preemp_1t_out		: OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
		tx_preemp_2t_out		: OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
		tx_vodctrl_out		: OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
	);
END reconfig_side;


ARCHITECTURE RTL OF reconfig_side IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "alt2gxb_reconfig";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "base_port_width=1;cbx_blackbox_list=-lpm_mux;channel_address_width=8;enable_chl_addr_for_analog_ctrl=TRUE;enable_dfe=ON;enable_eye_monitor=ON;enable_illegal_mode_check=TRUE;enable_self_recovery=TRUE;intended_device_family=Stratix IV;number_of_channels=144;number_of_reconfig_ports=36;read_base_port_width=1;reconfig_mode_sel_width=4;rx_eqdcgain_port_width=3;tx_preemp_port_width=5;enable_buf_cal=true;reconfig_fromgxb_width=612;reconfig_togxb_width=4;";
	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (4 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (2 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC ;
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (15 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC ;
	SIGNAL sub_wire6	: STD_LOGIC ;
	SIGNAL sub_wire7	: STD_LOGIC ;
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (4 DOWNTO 0);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (2 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (4 DOWNTO 0);



	COMPONENT reconfig_side_alt2gxb_reconfig_4og2
	PORT (
			ctrl_read	: IN STD_LOGIC ;
			logical_channel_address	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			reconfig_togxb	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			tx_preemp_1t	: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
			tx_preemp_2t_out	: OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
			tx_vodctrl_out	: OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			ctrl_writedata	: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			data_valid	: OUT STD_LOGIC ;
			reconfig_fromgxb	: IN STD_LOGIC_VECTOR (611 DOWNTO 0);
			tx_preemp_2t	: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
			tx_vodctrl	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			ctrl_address	: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
			ctrl_readdata	: OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			ctrl_waitrequest	: OUT STD_LOGIC ;
			error	: OUT STD_LOGIC ;
			busy	: OUT STD_LOGIC ;
			ctrl_write	: IN STD_LOGIC ;
			rx_eqctrl_out	: OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			tx_preemp_0t	: IN STD_LOGIC_VECTOR (4 DOWNTO 0);
			tx_preemp_1t_out	: OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
			write_all	: IN STD_LOGIC ;
			read	: IN STD_LOGIC ;
			reconfig_mode_sel	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			rx_eqctrl	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			rx_eqdcgain_out	: OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			rx_eqdcgain	: IN STD_LOGIC_VECTOR (2 DOWNTO 0);
			reconfig_clk	: IN STD_LOGIC ;
			tx_preemp_0t_out	: OUT STD_LOGIC_VECTOR (4 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	reconfig_togxb    <= sub_wire0(3 DOWNTO 0);
	tx_preemp_2t_out    <= sub_wire1(4 DOWNTO 0);
	tx_vodctrl_out    <= sub_wire2(2 DOWNTO 0);
	data_valid    <= sub_wire3;
	ctrl_readdata    <= sub_wire4(15 DOWNTO 0);
	ctrl_waitrequest    <= sub_wire5;
	error    <= sub_wire6;
	busy    <= sub_wire7;
	rx_eqctrl_out    <= sub_wire8(3 DOWNTO 0);
	tx_preemp_1t_out    <= sub_wire9(4 DOWNTO 0);
	rx_eqdcgain_out    <= sub_wire10(2 DOWNTO 0);
	tx_preemp_0t_out    <= sub_wire11(4 DOWNTO 0);

	reconfig_side_alt2gxb_reconfig_4og2_component : reconfig_side_alt2gxb_reconfig_4og2
	PORT MAP (
		ctrl_read => ctrl_read,
		logical_channel_address => logical_channel_address,
		tx_preemp_1t => tx_preemp_1t,
		ctrl_writedata => ctrl_writedata,
		reconfig_fromgxb => reconfig_fromgxb,
		tx_preemp_2t => tx_preemp_2t,
		tx_vodctrl => tx_vodctrl,
		ctrl_address => ctrl_address,
		ctrl_write => ctrl_write,
		tx_preemp_0t => tx_preemp_0t,
		write_all => write_all,
		read => read,
		reconfig_mode_sel => reconfig_mode_sel,
		rx_eqctrl => rx_eqctrl,
		rx_eqdcgain => rx_eqdcgain,
		reconfig_clk => reconfig_clk,
		reconfig_togxb => sub_wire0,
		tx_preemp_2t_out => sub_wire1,
		tx_vodctrl_out => sub_wire2,
		data_valid => sub_wire3,
		ctrl_readdata => sub_wire4,
		ctrl_waitrequest => sub_wire5,
		error => sub_wire6,
		busy => sub_wire7,
		rx_eqctrl_out => sub_wire8,
		tx_preemp_1t_out => sub_wire9,
		rx_eqdcgain_out => sub_wire10,
		tx_preemp_0t_out => sub_wire11
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: ADCE NUMERIC "0"
-- Retrieval info: PRIVATE: CMU_PLL NUMERIC "0"
-- Retrieval info: PRIVATE: DATA_RATE NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
-- Retrieval info: PRIVATE: PMA NUMERIC "1"
-- Retrieval info: PRIVATE: PROTO_SWITCH NUMERIC "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: CONSTANT: BASE_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: CBX_BLACKBOX_LIST STRING "-lpm_mux"
-- Retrieval info: CONSTANT: CHANNEL_ADDRESS_WIDTH NUMERIC "8"
-- Retrieval info: CONSTANT: ENABLE_CHL_ADDR_FOR_ANALOG_CTRL STRING "TRUE"
-- Retrieval info: CONSTANT: ENABLE_DFE STRING "ON"
-- Retrieval info: CONSTANT: ENABLE_EYE_MONITOR STRING "ON"
-- Retrieval info: CONSTANT: ENABLE_ILLEGAL_MODE_CHECK STRING "TRUE"
-- Retrieval info: CONSTANT: ENABLE_SELF_RECOVERY STRING "TRUE"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix IV"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "144"
-- Retrieval info: CONSTANT: NUMBER_OF_RECONFIG_PORTS NUMERIC "36"
-- Retrieval info: CONSTANT: READ_BASE_PORT_WIDTH NUMERIC "1"
-- Retrieval info: CONSTANT: RECONFIG_MODE_SEL_WIDTH NUMERIC "4"
-- Retrieval info: CONSTANT: RX_EQDCGAIN_PORT_WIDTH NUMERIC "3"
-- Retrieval info: CONSTANT: TX_PREEMP_PORT_WIDTH NUMERIC "5"
-- Retrieval info: CONSTANT: enable_buf_cal STRING "true"
-- Retrieval info: CONSTANT: reconfig_fromgxb_width NUMERIC "612"
-- Retrieval info: CONSTANT: reconfig_togxb_width NUMERIC "4"
-- Retrieval info: USED_PORT: busy 0 0 0 0 OUTPUT NODEFVAL "busy"
-- Retrieval info: USED_PORT: ctrl_address 0 0 16 0 INPUT NODEFVAL "ctrl_address[15..0]"
-- Retrieval info: USED_PORT: ctrl_read 0 0 0 0 INPUT NODEFVAL "ctrl_read"
-- Retrieval info: USED_PORT: ctrl_readdata 0 0 16 0 OUTPUT NODEFVAL "ctrl_readdata[15..0]"
-- Retrieval info: USED_PORT: ctrl_waitrequest 0 0 0 0 OUTPUT NODEFVAL "ctrl_waitrequest"
-- Retrieval info: USED_PORT: ctrl_write 0 0 0 0 INPUT NODEFVAL "ctrl_write"
-- Retrieval info: USED_PORT: ctrl_writedata 0 0 16 0 INPUT NODEFVAL "ctrl_writedata[15..0]"
-- Retrieval info: USED_PORT: data_valid 0 0 0 0 OUTPUT NODEFVAL "data_valid"
-- Retrieval info: USED_PORT: error 0 0 0 0 OUTPUT NODEFVAL "error"
-- Retrieval info: USED_PORT: logical_channel_address 0 0 8 0 INPUT NODEFVAL "logical_channel_address[7..0]"
-- Retrieval info: USED_PORT: read 0 0 0 0 INPUT NODEFVAL "read"
-- Retrieval info: USED_PORT: reconfig_clk 0 0 0 0 INPUT NODEFVAL "reconfig_clk"
-- Retrieval info: USED_PORT: reconfig_fromgxb 0 0 612 0 INPUT NODEFVAL "reconfig_fromgxb[611..0]"
-- Retrieval info: USED_PORT: reconfig_mode_sel 0 0 4 0 INPUT NODEFVAL "reconfig_mode_sel[3..0]"
-- Retrieval info: USED_PORT: reconfig_togxb 0 0 4 0 OUTPUT NODEFVAL "reconfig_togxb[3..0]"
-- Retrieval info: USED_PORT: rx_eqctrl 0 0 4 0 INPUT NODEFVAL "rx_eqctrl[3..0]"
-- Retrieval info: USED_PORT: rx_eqctrl_out 0 0 4 0 OUTPUT NODEFVAL "rx_eqctrl_out[3..0]"
-- Retrieval info: USED_PORT: rx_eqdcgain 0 0 3 0 INPUT NODEFVAL "rx_eqdcgain[2..0]"
-- Retrieval info: USED_PORT: rx_eqdcgain_out 0 0 3 0 OUTPUT NODEFVAL "rx_eqdcgain_out[2..0]"
-- Retrieval info: USED_PORT: tx_preemp_0t 0 0 5 0 INPUT NODEFVAL "tx_preemp_0t[4..0]"
-- Retrieval info: USED_PORT: tx_preemp_0t_out 0 0 5 0 OUTPUT NODEFVAL "tx_preemp_0t_out[4..0]"
-- Retrieval info: USED_PORT: tx_preemp_1t 0 0 5 0 INPUT NODEFVAL "tx_preemp_1t[4..0]"
-- Retrieval info: USED_PORT: tx_preemp_1t_out 0 0 5 0 OUTPUT NODEFVAL "tx_preemp_1t_out[4..0]"
-- Retrieval info: USED_PORT: tx_preemp_2t 0 0 5 0 INPUT NODEFVAL "tx_preemp_2t[4..0]"
-- Retrieval info: USED_PORT: tx_preemp_2t_out 0 0 5 0 OUTPUT NODEFVAL "tx_preemp_2t_out[4..0]"
-- Retrieval info: USED_PORT: tx_vodctrl 0 0 3 0 INPUT NODEFVAL "tx_vodctrl[2..0]"
-- Retrieval info: USED_PORT: tx_vodctrl_out 0 0 3 0 OUTPUT NODEFVAL "tx_vodctrl_out[2..0]"
-- Retrieval info: USED_PORT: write_all 0 0 0 0 INPUT NODEFVAL "write_all"
-- Retrieval info: CONNECT: @ctrl_address 0 0 16 0 ctrl_address 0 0 16 0
-- Retrieval info: CONNECT: @ctrl_read 0 0 0 0 ctrl_read 0 0 0 0
-- Retrieval info: CONNECT: @ctrl_write 0 0 0 0 ctrl_write 0 0 0 0
-- Retrieval info: CONNECT: @ctrl_writedata 0 0 16 0 ctrl_writedata 0 0 16 0
-- Retrieval info: CONNECT: @logical_channel_address 0 0 8 0 logical_channel_address 0 0 8 0
-- Retrieval info: CONNECT: @read 0 0 0 0 read 0 0 0 0
-- Retrieval info: CONNECT: @reconfig_clk 0 0 0 0 reconfig_clk 0 0 0 0
-- Retrieval info: CONNECT: @reconfig_fromgxb 0 0 612 0 reconfig_fromgxb 0 0 612 0
-- Retrieval info: CONNECT: @reconfig_mode_sel 0 0 4 0 reconfig_mode_sel 0 0 4 0
-- Retrieval info: CONNECT: @rx_eqctrl 0 0 4 0 rx_eqctrl 0 0 4 0
-- Retrieval info: CONNECT: @rx_eqdcgain 0 0 3 0 rx_eqdcgain 0 0 3 0
-- Retrieval info: CONNECT: @tx_preemp_0t 0 0 5 0 tx_preemp_0t 0 0 5 0
-- Retrieval info: CONNECT: @tx_preemp_1t 0 0 5 0 tx_preemp_1t 0 0 5 0
-- Retrieval info: CONNECT: @tx_preemp_2t 0 0 5 0 tx_preemp_2t 0 0 5 0
-- Retrieval info: CONNECT: @tx_vodctrl 0 0 3 0 tx_vodctrl 0 0 3 0
-- Retrieval info: CONNECT: @write_all 0 0 0 0 write_all 0 0 0 0
-- Retrieval info: CONNECT: busy 0 0 0 0 @busy 0 0 0 0
-- Retrieval info: CONNECT: ctrl_readdata 0 0 16 0 @ctrl_readdata 0 0 16 0
-- Retrieval info: CONNECT: ctrl_waitrequest 0 0 0 0 @ctrl_waitrequest 0 0 0 0
-- Retrieval info: CONNECT: data_valid 0 0 0 0 @data_valid 0 0 0 0
-- Retrieval info: CONNECT: error 0 0 0 0 @error 0 0 0 0
-- Retrieval info: CONNECT: reconfig_togxb 0 0 4 0 @reconfig_togxb 0 0 4 0
-- Retrieval info: CONNECT: rx_eqctrl_out 0 0 4 0 @rx_eqctrl_out 0 0 4 0
-- Retrieval info: CONNECT: rx_eqdcgain_out 0 0 3 0 @rx_eqdcgain_out 0 0 3 0
-- Retrieval info: CONNECT: tx_preemp_0t_out 0 0 5 0 @tx_preemp_0t_out 0 0 5 0
-- Retrieval info: CONNECT: tx_preemp_1t_out 0 0 5 0 @tx_preemp_1t_out 0 0 5 0
-- Retrieval info: CONNECT: tx_preemp_2t_out 0 0 5 0 @tx_preemp_2t_out 0 0 5 0
-- Retrieval info: CONNECT: tx_vodctrl_out 0 0 3 0 @tx_vodctrl_out 0 0 3 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL reconfig_side.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL reconfig_side.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL reconfig_side.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL reconfig_side.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL reconfig_side_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
-- Retrieval info: LIB_FILE: lpm
