-- sopc_system.vhd

-- Generated using ACDS version 13.0sp1 232 at 2015.06.12.15:50:13

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sopc_system is
	port (
		clk_in_reset_reset_n            : in    std_logic                     := '0';             -- clk_in_reset.reset_n
		clk_in_clk                      : in    std_logic                     := '0';             --       clk_in.clk
		ddr2_status_local_init_done     : out   std_logic;                                        --  ddr2_status.local_init_done
		ddr2_status_local_cal_success   : out   std_logic;                                        --             .local_cal_success
		ddr2_status_local_cal_fail      : out   std_logic;                                        --             .local_cal_fail
		ddr2_mem_mem_a                  : out   std_logic_vector(12 downto 0);                    --     ddr2_mem.mem_a
		ddr2_mem_mem_ba                 : out   std_logic_vector(2 downto 0);                     --             .mem_ba
		ddr2_mem_mem_ck                 : out   std_logic_vector(0 downto 0);                     --             .mem_ck
		ddr2_mem_mem_ck_n               : out   std_logic_vector(0 downto 0);                     --             .mem_ck_n
		ddr2_mem_mem_cke                : out   std_logic_vector(0 downto 0);                     --             .mem_cke
		ddr2_mem_mem_cs_n               : out   std_logic_vector(0 downto 0);                     --             .mem_cs_n
		ddr2_mem_mem_dm                 : out   std_logic_vector(1 downto 0);                     --             .mem_dm
		ddr2_mem_mem_ras_n              : out   std_logic_vector(0 downto 0);                     --             .mem_ras_n
		ddr2_mem_mem_cas_n              : out   std_logic_vector(0 downto 0);                     --             .mem_cas_n
		ddr2_mem_mem_we_n               : out   std_logic_vector(0 downto 0);                     --             .mem_we_n
		ddr2_mem_mem_dq                 : inout std_logic_vector(15 downto 0) := (others => '0'); --             .mem_dq
		ddr2_mem_mem_dqs                : inout std_logic_vector(1 downto 0)  := (others => '0'); --             .mem_dqs
		ddr2_mem_mem_dqs_n              : inout std_logic_vector(1 downto 0)  := (others => '0'); --             .mem_dqs_n
		ddr2_mem_mem_odt                : out   std_logic_vector(0 downto 0);                     --             .mem_odt
		cfi_tcm_address_out             : out   std_logic_vector(26 downto 0);                    --          cfi.tcm_address_out
		cfi_tcm_outputenable_n_out      : out   std_logic_vector(0 downto 0);                     --             .tcm_outputenable_n_out
		cfi_tcm_reset_n_out             : out   std_logic_vector(0 downto 0);                     --             .tcm_reset_n_out
		cfi_tcm_write_n_out             : out   std_logic_vector(0 downto 0);                     --             .tcm_write_n_out
		cfi_tcm_data_out                : inout std_logic_vector(15 downto 0) := (others => '0'); --             .tcm_data_out
		cfi_tcm_chipselect_n_out        : out   std_logic_vector(0 downto 0);                     --             .tcm_chipselect_n_out
		ddr2_oct_rdn                    : in    std_logic                     := '0';             --     ddr2_oct.rdn
		ddr2_oct_rup                    : in    std_logic                     := '0';             --             .rup
		gtpbus_CLK                      : out   std_logic;                                        --       gtpbus.CLK
		gtpbus_RESET                    : out   std_logic;                                        --             .RESET
		gtpbus_DIN                      : out   std_logic_vector(31 downto 0);                    --             .DIN
		gtpbus_DOUT                     : in    std_logic_vector(31 downto 0) := (others => '0'); --             .DOUT
		gtpbus_WR                       : out   std_logic;                                        --             .WR
		gtpbus_RD                       : out   std_logic;                                        --             .RD
		gtpbus_ACK                      : in    std_logic                     := '0';             --             .ACK
		gtpbus_ADDR                     : out   std_logic_vector(15 downto 0);                    --             .ADDR
		gtpbus_IRQ                      : in    std_logic                     := '0';             --             .IRQ
		tse_mdio_mdc                    : out   std_logic;                                        --     tse_mdio.mdc
		tse_mdio_mdio_in                : in    std_logic                     := '0';             --             .mdio_in
		tse_mdio_mdio_out               : out   std_logic;                                        --             .mdio_out
		tse_mdio_mdio_oen               : out   std_logic;                                        --             .mdio_oen
		tse_rgmii_rgmii_in              : in    std_logic_vector(3 downto 0)  := (others => '0'); --    tse_rgmii.rgmii_in
		tse_rgmii_rgmii_out             : out   std_logic_vector(3 downto 0);                     --             .rgmii_out
		tse_rgmii_rx_control            : in    std_logic                     := '0';             --             .rx_control
		tse_rgmii_tx_control            : out   std_logic;                                        --             .tx_control
		tse_status_set_10               : in    std_logic                     := '0';             --   tse_status.set_10
		tse_status_set_1000             : in    std_logic                     := '0';             --             .set_1000
		tse_status_eth_mode             : out   std_logic;                                        --             .eth_mode
		tse_status_ena_10               : out   std_logic;                                        --             .ena_10
		tse_txclk_clk                   : in    std_logic                     := '0';             --    tse_txclk.clk
		tse_rxclk_clk                   : in    std_logic                     := '0';             --    tse_rxclk.clk
		cfi_fpga_tcm_address_out        : out   std_logic_vector(26 downto 0);                    --     cfi_fpga.tcm_address_out
		cfi_fpga_tcm_outputenable_n_out : out   std_logic_vector(0 downto 0);                     --             .tcm_outputenable_n_out
		cfi_fpga_tcm_reset_n_out        : out   std_logic_vector(0 downto 0);                     --             .tcm_reset_n_out
		cfi_fpga_tcm_write_n_out        : out   std_logic_vector(0 downto 0);                     --             .tcm_write_n_out
		cfi_fpga_tcm_data_out           : inout std_logic_vector(15 downto 0) := (others => '0'); --             .tcm_data_out
		cfi_fpga_tcm_chipselect_n_out   : out   std_logic_vector(0 downto 0);                     --             .tcm_chipselect_n_out
		tse_misc_xon_gen                : in    std_logic                     := '0';             --     tse_misc.xon_gen
		tse_misc_xoff_gen               : in    std_logic                     := '0';             --             .xoff_gen
		tse_misc_magic_wakeup           : out   std_logic;                                        --             .magic_wakeup
		tse_misc_magic_sleep_n          : in    std_logic                     := '0';             --             .magic_sleep_n
		tse_misc_ff_tx_crc_fwd          : in    std_logic                     := '0';             --             .ff_tx_crc_fwd
		tse_misc_ff_tx_septy            : out   std_logic;                                        --             .ff_tx_septy
		tse_misc_tx_ff_uflow            : out   std_logic;                                        --             .tx_ff_uflow
		tse_misc_ff_tx_a_full           : out   std_logic;                                        --             .ff_tx_a_full
		tse_misc_ff_tx_a_empty          : out   std_logic;                                        --             .ff_tx_a_empty
		tse_misc_rx_err_stat            : out   std_logic_vector(17 downto 0);                    --             .rx_err_stat
		tse_misc_rx_frm_type            : out   std_logic_vector(3 downto 0);                     --             .rx_frm_type
		tse_misc_ff_rx_dsav             : out   std_logic;                                        --             .ff_rx_dsav
		tse_misc_ff_rx_a_full           : out   std_logic;                                        --             .ff_rx_a_full
		tse_misc_ff_rx_a_empty          : out   std_logic                                         --             .ff_rx_a_empty
	);
end entity sopc_system;

architecture rtl of sopc_system is
	component sopc_system_linux_timer_1ms is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component sopc_system_linux_timer_1ms;

	component sopc_system_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component sopc_system_jtag_uart;

	component sopc_system_sgdma_rx is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			in_startofpacket              : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket                : in  std_logic                     := 'X';             -- endofpacket
			in_data                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_valid                      : in  std_logic                     := 'X';             -- valid
			in_ready                      : out std_logic;                                        -- ready
			in_empty                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			in_error                      : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- error
			m_write_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			m_write_address               : out std_logic_vector(31 downto 0);                    -- address
			m_write_write                 : out std_logic;                                        -- write
			m_write_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			m_write_byteenable            : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component sopc_system_sgdma_rx;

	component sopc_system_sgdma_tx is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			m_read_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m_read_readdatavalid          : in  std_logic                     := 'X';             -- readdatavalid
			m_read_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			m_read_address                : out std_logic_vector(31 downto 0);                    -- address
			m_read_read                   : out std_logic;                                        -- read
			out_data                      : out std_logic_vector(31 downto 0);                    -- data
			out_valid                     : out std_logic;                                        -- valid
			out_ready                     : in  std_logic                     := 'X';             -- ready
			out_endofpacket               : out std_logic;                                        -- endofpacket
			out_startofpacket             : out std_logic;                                        -- startofpacket
			out_empty                     : out std_logic_vector(1 downto 0);                     -- empty
			out_error                     : out std_logic                                         -- error
		);
	end component sopc_system_sgdma_tx;

	component sopc_system_descriptor_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component sopc_system_descriptor_memory;

	component sopc_system_linux_cpu is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(28 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(28 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			dcm0_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			dcm0_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			dcm0_readdatavalid                    : in  std_logic                     := 'X';             -- readdatavalid
			dcm0_address                          : out std_logic_vector(28 downto 0);                    -- address
			dcm0_read                             : out std_logic;                                        -- read
			dcm0_clken                            : out std_logic;                                        -- clken
			dcm0_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			dcm0_write                            : out std_logic;                                        -- write
			dcm0_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			icm0_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			icm0_waitrequest                      : in  std_logic                     := 'X';             -- waitrequest
			icm0_readdatavalid                    : in  std_logic                     := 'X';             -- readdatavalid
			icm0_address                          : out std_logic_vector(28 downto 0);                    -- address
			icm0_read                             : out std_logic;                                        -- read
			icm0_clken                            : out std_logic;                                        -- clken
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component sopc_system_linux_cpu;

	component sopc_system_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component sopc_system_sysid;

	component sopc_system_sdram_0 is
		port (
			pll_ref_clk        : in    std_logic                     := 'X';             -- clk
			global_reset_n     : in    std_logic                     := 'X';             -- reset_n
			soft_reset_n       : in    std_logic                     := 'X';             -- reset_n
			afi_clk            : out   std_logic;                                        -- clk
			afi_half_clk       : out   std_logic;                                        -- clk
			afi_reset_n        : out   std_logic;                                        -- reset_n
			afi_reset_export_n : out   std_logic;                                        -- reset_n
			mem_a              : out   std_logic_vector(12 downto 0);                    -- mem_a
			mem_ba             : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck             : out   std_logic_vector(0 downto 0);                     -- mem_ck
			mem_ck_n           : out   std_logic_vector(0 downto 0);                     -- mem_ck_n
			mem_cke            : out   std_logic_vector(0 downto 0);                     -- mem_cke
			mem_cs_n           : out   std_logic_vector(0 downto 0);                     -- mem_cs_n
			mem_dm             : out   std_logic_vector(1 downto 0);                     -- mem_dm
			mem_ras_n          : out   std_logic_vector(0 downto 0);                     -- mem_ras_n
			mem_cas_n          : out   std_logic_vector(0 downto 0);                     -- mem_cas_n
			mem_we_n           : out   std_logic_vector(0 downto 0);                     -- mem_we_n
			mem_dq             : inout std_logic_vector(15 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs            : inout std_logic_vector(1 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n          : inout std_logic_vector(1 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt            : out   std_logic_vector(0 downto 0);                     -- mem_odt
			avl_ready          : out   std_logic;                                        -- waitrequest_n
			avl_burstbegin     : in    std_logic                     := 'X';             -- beginbursttransfer
			avl_addr           : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			avl_rdata_valid    : out   std_logic;                                        -- readdatavalid
			avl_rdata          : out   std_logic_vector(63 downto 0);                    -- readdata
			avl_wdata          : in    std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			avl_be             : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req       : in    std_logic                     := 'X';             -- read
			avl_write_req      : in    std_logic                     := 'X';             -- write
			avl_size           : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			local_init_done    : out   std_logic;                                        -- local_init_done
			local_cal_success  : out   std_logic;                                        -- local_cal_success
			local_cal_fail     : out   std_logic;                                        -- local_cal_fail
			oct_rdn            : in    std_logic                     := 'X';             -- rdn
			oct_rup            : in    std_logic                     := 'X'              -- rup
		);
	end component sopc_system_sdram_0;

	component sopc_system_cfi_flash_ts_controller is
		generic (
			TCM_ADDRESS_W                  : integer := 30;
			TCM_DATA_W                     : integer := 32;
			TCM_BYTEENABLE_W               : integer := 4;
			TCM_READ_WAIT                  : integer := 1;
			TCM_WRITE_WAIT                 : integer := 0;
			TCM_SETUP_WAIT                 : integer := 0;
			TCM_DATA_HOLD                  : integer := 0;
			TCM_TURNAROUND_TIME            : integer := 2;
			TCM_TIMING_UNITS               : integer := 1;
			TCM_READLATENCY                : integer := 2;
			TCM_SYMBOLS_PER_WORD           : integer := 4;
			USE_READDATA                   : integer := 1;
			USE_WRITEDATA                  : integer := 1;
			USE_READ                       : integer := 1;
			USE_WRITE                      : integer := 1;
			USE_BYTEENABLE                 : integer := 1;
			USE_CHIPSELECT                 : integer := 0;
			USE_LOCK                       : integer := 0;
			USE_ADDRESS                    : integer := 1;
			USE_WAITREQUEST                : integer := 0;
			USE_WRITEBYTEENABLE            : integer := 0;
			USE_OUTPUTENABLE               : integer := 0;
			USE_RESETREQUEST               : integer := 0;
			USE_IRQ                        : integer := 0;
			USE_RESET_OUTPUT               : integer := 0;
			ACTIVE_LOW_READ                : integer := 0;
			ACTIVE_LOW_LOCK                : integer := 0;
			ACTIVE_LOW_WRITE               : integer := 0;
			ACTIVE_LOW_CHIPSELECT          : integer := 0;
			ACTIVE_LOW_BYTEENABLE          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE        : integer := 0;
			ACTIVE_LOW_WRITEBYTEENABLE     : integer := 0;
			ACTIVE_LOW_WAITREQUEST         : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER       : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0
		);
		port (
			clk_clk                : in  std_logic                     := 'X';             -- clk
			reset_reset            : in  std_logic                     := 'X';             -- reset
			uas_address            : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			uas_burstcount         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uas_read               : in  std_logic                     := 'X';             -- read
			uas_write              : in  std_logic                     := 'X';             -- write
			uas_waitrequest        : out std_logic;                                        -- waitrequest
			uas_readdatavalid      : out std_logic;                                        -- readdatavalid
			uas_byteenable         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uas_readdata           : out std_logic_vector(15 downto 0);                    -- readdata
			uas_writedata          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uas_lock               : in  std_logic                     := 'X';             -- lock
			uas_debugaccess        : in  std_logic                     := 'X';             -- debugaccess
			tcm_write_n_out        : out std_logic;                                        -- write_n_out
			tcm_chipselect_n_out   : out std_logic;                                        -- chipselect_n_out
			tcm_outputenable_n_out : out std_logic;                                        -- outputenable_n_out
			tcm_reset_n_out        : out std_logic;                                        -- reset_n_out
			tcm_request            : out std_logic;                                        -- request
			tcm_grant              : in  std_logic                     := 'X';             -- grant
			tcm_address_out        : out std_logic_vector(26 downto 0);                    -- address_out
			tcm_data_out           : out std_logic_vector(15 downto 0);                    -- data_out
			tcm_data_outen         : out std_logic;                                        -- data_outen
			tcm_data_in            : in  std_logic_vector(15 downto 0) := (others => 'X')  -- data_in
		);
	end component sopc_system_cfi_flash_ts_controller;

	component sopc_system_cfi_flash_ts_bridge is
		port (
			clk                        : in    std_logic                     := 'X';             -- clk
			reset                      : in    std_logic                     := 'X';             -- reset
			request                    : in    std_logic                     := 'X';             -- request
			grant                      : out   std_logic;                                        -- grant
			tcs_tcm_address_out        : in    std_logic_vector(26 downto 0) := (others => 'X'); -- address_out
			tcs_tcm_outputenable_n_out : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- outputenable_n_out
			tcs_tcm_reset_n_out        : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- reset_n_out
			tcs_tcm_write_n_out        : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_out
			tcs_tcm_data_out           : in    std_logic_vector(15 downto 0) := (others => 'X'); -- data_out
			tcs_tcm_data_outen         : in    std_logic                     := 'X';             -- data_outen
			tcs_tcm_data_in            : out   std_logic_vector(15 downto 0);                    -- data_in
			tcs_tcm_chipselect_n_out   : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- chipselect_n_out
			tcm_address_out            : out   std_logic_vector(26 downto 0);                    -- tcm_address_out
			tcm_outputenable_n_out     : out   std_logic_vector(0 downto 0);                     -- tcm_outputenable_n_out
			tcm_reset_n_out            : out   std_logic_vector(0 downto 0);                     -- tcm_reset_n_out
			tcm_write_n_out            : out   std_logic_vector(0 downto 0);                     -- tcm_write_n_out
			tcm_data_out               : inout std_logic_vector(15 downto 0) := (others => 'X'); -- tcm_data_out
			tcm_chipselect_n_out       : out   std_logic_vector(0 downto 0)                      -- tcm_chipselect_n_out
		);
	end component sopc_system_cfi_flash_ts_bridge;

	component gtp_regif is
		port (
			avs_s0_address     : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			avs_s0_read        : in  std_logic                     := 'X';             -- read
			avs_s0_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			avs_s0_write       : in  std_logic                     := 'X';             -- write
			avs_s0_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_s0_waitrequest : out std_logic;                                        -- waitrequest
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			BUS_CLK            : out std_logic;                                        -- export
			BUS_RESET          : out std_logic;                                        -- export
			BUS_DIN            : out std_logic_vector(31 downto 0);                    -- export
			BUS_DOUT           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- export
			BUS_WR             : out std_logic;                                        -- export
			BUS_RD             : out std_logic;                                        -- export
			BUS_ACK            : in  std_logic                     := 'X';             -- export
			BUS_ADDR           : out std_logic_vector(15 downto 0);                    -- export
			BUS_IRQ            : in  std_logic                     := 'X';             -- export
			irq                : out std_logic                                         -- irq
		);
	end component gtp_regif;

	component sopc_system_tse_mac is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			address       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			read          : in  std_logic                     := 'X';             -- read
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			write         : in  std_logic                     := 'X';             -- write
			waitrequest   : out std_logic;                                        -- waitrequest
			tx_clk        : in  std_logic                     := 'X';             -- clk
			rx_clk        : in  std_logic                     := 'X';             -- clk
			set_10        : in  std_logic                     := 'X';             -- set_10
			set_1000      : in  std_logic                     := 'X';             -- set_1000
			eth_mode      : out std_logic;                                        -- eth_mode
			ena_10        : out std_logic;                                        -- ena_10
			rgmii_in      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- rgmii_in
			rgmii_out     : out std_logic_vector(3 downto 0);                     -- rgmii_out
			rx_control    : in  std_logic                     := 'X';             -- rx_control
			tx_control    : out std_logic;                                        -- tx_control
			ff_rx_clk     : in  std_logic                     := 'X';             -- clk
			ff_tx_clk     : in  std_logic                     := 'X';             -- clk
			ff_rx_data    : out std_logic_vector(31 downto 0);                    -- data
			ff_rx_eop     : out std_logic;                                        -- endofpacket
			rx_err        : out std_logic_vector(5 downto 0);                     -- error
			ff_rx_mod     : out std_logic_vector(1 downto 0);                     -- empty
			ff_rx_rdy     : in  std_logic                     := 'X';             -- ready
			ff_rx_sop     : out std_logic;                                        -- startofpacket
			ff_rx_dval    : out std_logic;                                        -- valid
			ff_tx_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			ff_tx_eop     : in  std_logic                     := 'X';             -- endofpacket
			ff_tx_err     : in  std_logic                     := 'X';             -- error
			ff_tx_mod     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			ff_tx_rdy     : out std_logic;                                        -- ready
			ff_tx_sop     : in  std_logic                     := 'X';             -- startofpacket
			ff_tx_wren    : in  std_logic                     := 'X';             -- valid
			mdc           : out std_logic;                                        -- mdc
			mdio_in       : in  std_logic                     := 'X';             -- mdio_in
			mdio_out      : out std_logic;                                        -- mdio_out
			mdio_oen      : out std_logic;                                        -- mdio_oen
			xon_gen       : in  std_logic                     := 'X';             -- xon_gen
			xoff_gen      : in  std_logic                     := 'X';             -- xoff_gen
			magic_wakeup  : out std_logic;                                        -- magic_wakeup
			magic_sleep_n : in  std_logic                     := 'X';             -- magic_sleep_n
			ff_tx_crc_fwd : in  std_logic                     := 'X';             -- ff_tx_crc_fwd
			ff_tx_septy   : out std_logic;                                        -- ff_tx_septy
			tx_ff_uflow   : out std_logic;                                        -- tx_ff_uflow
			ff_tx_a_full  : out std_logic;                                        -- ff_tx_a_full
			ff_tx_a_empty : out std_logic;                                        -- ff_tx_a_empty
			rx_err_stat   : out std_logic_vector(17 downto 0);                    -- rx_err_stat
			rx_frm_type   : out std_logic_vector(3 downto 0);                     -- rx_frm_type
			ff_rx_dsav    : out std_logic;                                        -- ff_rx_dsav
			ff_rx_a_full  : out std_logic;                                        -- ff_rx_a_full
			ff_rx_a_empty : out std_logic                                         -- ff_rx_a_empty
		);
	end component sopc_system_tse_mac;

	component sopc_system_cfi_flash_ts_bridge_fpga is
		port (
			clk                        : in    std_logic                     := 'X';             -- clk
			reset                      : in    std_logic                     := 'X';             -- reset
			request                    : in    std_logic                     := 'X';             -- request
			grant                      : out   std_logic;                                        -- grant
			tcs_tcm_address_out        : in    std_logic_vector(26 downto 0) := (others => 'X'); -- address_out
			tcs_tcm_outputenable_n_out : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- outputenable_n_out
			tcs_tcm_reset_n_out        : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- reset_n_out
			tcs_tcm_write_n_out        : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_out
			tcs_tcm_data_out           : in    std_logic_vector(15 downto 0) := (others => 'X'); -- data_out
			tcs_tcm_data_outen         : in    std_logic                     := 'X';             -- data_outen
			tcs_tcm_data_in            : out   std_logic_vector(15 downto 0);                    -- data_in
			tcs_tcm_chipselect_n_out   : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- chipselect_n_out
			tcm_address_out            : out   std_logic_vector(26 downto 0);                    -- tcm_address_out
			tcm_outputenable_n_out     : out   std_logic_vector(0 downto 0);                     -- tcm_outputenable_n_out
			tcm_reset_n_out            : out   std_logic_vector(0 downto 0);                     -- tcm_reset_n_out
			tcm_write_n_out            : out   std_logic_vector(0 downto 0);                     -- tcm_write_n_out
			tcm_data_out               : inout std_logic_vector(15 downto 0) := (others => 'X'); -- tcm_data_out
			tcm_chipselect_n_out       : out   std_logic_vector(0 downto 0)                      -- tcm_chipselect_n_out
		);
	end component sopc_system_cfi_flash_ts_bridge_fpga;

	component sopc_system_tlb_miss_ram_1k is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X'              -- reset_req
		);
	end component sopc_system_tlb_miss_ram_1k;

	component sopc_system_addr_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(99 downto 0);                    -- data
			src_channel        : out std_logic_vector(3 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component sopc_system_addr_router;

	component sopc_system_addr_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(99 downto 0);                    -- data
			src_channel        : out std_logic_vector(3 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component sopc_system_addr_router_001;

	component sopc_system_id_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(99 downto 0);                    -- data
			src_channel        : out std_logic_vector(3 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component sopc_system_id_router;

	component sopc_system_id_router_002 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(99 downto 0);                    -- data
			src_channel        : out std_logic_vector(3 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component sopc_system_id_router_002;

	component sopc_system_addr_router_002 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(100 downto 0);                    -- data
			src_channel        : out std_logic_vector(3 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component sopc_system_addr_router_002;

	component sopc_system_id_router_004 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(100 downto 0);                    -- data
			src_channel        : out std_logic_vector(3 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component sopc_system_id_router_004;

	component sopc_system_addr_router_006 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(93 downto 0);                    -- data
			src_channel        : out std_logic_vector(7 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component sopc_system_addr_router_006;

	component sopc_system_addr_router_007 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(93 downto 0);                    -- data
			src_channel        : out std_logic_vector(7 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component sopc_system_addr_router_007;

	component sopc_system_id_router_005 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(93 downto 0);                    -- data
			src_channel        : out std_logic_vector(7 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component sopc_system_id_router_005;

	component sopc_system_id_router_006 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(93 downto 0);                    -- data
			src_channel        : out std_logic_vector(7 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component sopc_system_id_router_006;

	component sopc_system_addr_router_008 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(94 downto 0);                    -- data
			src_channel        : out std_logic_vector(1 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component sopc_system_addr_router_008;

	component sopc_system_id_router_013 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(76 downto 0);                    -- data
			src_channel        : out std_logic_vector(1 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component sopc_system_id_router_013;

	component sopc_system_addr_router_009 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(98 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(98 downto 0);                    -- data
			src_channel        : out std_logic_vector(1 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component sopc_system_addr_router_009;

	component sopc_system_id_router_015 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(98 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(98 downto 0);                    -- data
			src_channel        : out std_logic_vector(1 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component sopc_system_id_router_015;

	component sopc_system_addr_router_011 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(96 downto 0);                    -- data
			src_channel        : out std_logic_vector(1 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component sopc_system_addr_router_011;

	component sopc_system_id_router_016 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(132 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(132 downto 0);                    -- data
			src_channel        : out std_logic_vector(1 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component sopc_system_id_router_016;

	component altera_merlin_burst_adapter is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(76 downto 0);                    -- data
			source0_channel       : out std_logic_vector(1 downto 0);                     -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component altera_merlin_burst_adapter;

	component sopc_system_cmd_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- data
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(99 downto 0);                    -- data
			src0_channel       : out std_logic_vector(3 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(99 downto 0);                    -- data
			src1_channel       : out std_logic_vector(3 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic;                                        -- endofpacket
			src2_ready         : in  std_logic                     := 'X';             -- ready
			src2_valid         : out std_logic;                                        -- valid
			src2_data          : out std_logic_vector(99 downto 0);                    -- data
			src2_channel       : out std_logic_vector(3 downto 0);                     -- channel
			src2_startofpacket : out std_logic;                                        -- startofpacket
			src2_endofpacket   : out std_logic;                                        -- endofpacket
			src3_ready         : in  std_logic                     := 'X';             -- ready
			src3_valid         : out std_logic;                                        -- valid
			src3_data          : out std_logic_vector(99 downto 0);                    -- data
			src3_channel       : out std_logic_vector(3 downto 0);                     -- channel
			src3_startofpacket : out std_logic;                                        -- startofpacket
			src3_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component sopc_system_cmd_xbar_demux;

	component sopc_system_cmd_xbar_demux_001 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- data
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(99 downto 0);                    -- data
			src0_channel       : out std_logic_vector(3 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(99 downto 0);                    -- data
			src1_channel       : out std_logic_vector(3 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic;                                        -- endofpacket
			src2_ready         : in  std_logic                     := 'X';             -- ready
			src2_valid         : out std_logic;                                        -- valid
			src2_data          : out std_logic_vector(99 downto 0);                    -- data
			src2_channel       : out std_logic_vector(3 downto 0);                     -- channel
			src2_startofpacket : out std_logic;                                        -- startofpacket
			src2_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component sopc_system_cmd_xbar_demux_001;

	component sopc_system_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(99 downto 0);                    -- data
			src_channel         : out std_logic_vector(3 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component sopc_system_cmd_xbar_mux;

	component sopc_system_rsp_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(99 downto 0);                    -- data
			src0_channel       : out std_logic_vector(3 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(99 downto 0);                    -- data
			src1_channel       : out std_logic_vector(3 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component sopc_system_rsp_xbar_demux;

	component sopc_system_rsp_xbar_demux_002 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(99 downto 0);                    -- data
			src0_channel       : out std_logic_vector(3 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component sopc_system_rsp_xbar_demux_002;

	component sopc_system_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(99 downto 0);                    -- data
			src_channel         : out std_logic_vector(3 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                        -- ready
			sink2_valid         : in  std_logic                     := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                        -- ready
			sink3_valid         : in  std_logic                     := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component sopc_system_rsp_xbar_mux;

	component sopc_system_rsp_xbar_mux_001 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(99 downto 0);                    -- data
			src_channel         : out std_logic_vector(3 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                        -- ready
			sink2_valid         : in  std_logic                     := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component sopc_system_rsp_xbar_mux_001;

	component sopc_system_cmd_xbar_demux_002 is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(100 downto 0);                    -- data
			src0_channel       : out std_logic_vector(3 downto 0);                      -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component sopc_system_cmd_xbar_demux_002;

	component sopc_system_cmd_xbar_mux_004 is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(100 downto 0);                    -- data
			src_channel         : out std_logic_vector(3 downto 0);                      -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                         -- ready
			sink2_valid         : in  std_logic                      := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                         -- ready
			sink3_valid         : in  std_logic                      := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component sopc_system_cmd_xbar_mux_004;

	component sopc_system_rsp_xbar_demux_004 is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(100 downto 0);                    -- data
			src0_channel       : out std_logic_vector(3 downto 0);                      -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(100 downto 0);                    -- data
			src1_channel       : out std_logic_vector(3 downto 0);                      -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic;                                         -- endofpacket
			src2_ready         : in  std_logic                      := 'X';             -- ready
			src2_valid         : out std_logic;                                         -- valid
			src2_data          : out std_logic_vector(100 downto 0);                    -- data
			src2_channel       : out std_logic_vector(3 downto 0);                      -- channel
			src2_startofpacket : out std_logic;                                         -- startofpacket
			src2_endofpacket   : out std_logic;                                         -- endofpacket
			src3_ready         : in  std_logic                      := 'X';             -- ready
			src3_valid         : out std_logic;                                         -- valid
			src3_data          : out std_logic_vector(100 downto 0);                    -- data
			src3_channel       : out std_logic_vector(3 downto 0);                      -- channel
			src3_startofpacket : out std_logic;                                         -- startofpacket
			src3_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component sopc_system_rsp_xbar_demux_004;

	component sopc_system_cmd_xbar_demux_006 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(93 downto 0);                    -- data
			src0_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component sopc_system_cmd_xbar_demux_006;

	component sopc_system_cmd_xbar_demux_007 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(93 downto 0);                    -- data
			src0_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(93 downto 0);                    -- data
			src1_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic;                                        -- endofpacket
			src2_ready         : in  std_logic                     := 'X';             -- ready
			src2_valid         : out std_logic;                                        -- valid
			src2_data          : out std_logic_vector(93 downto 0);                    -- data
			src2_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src2_startofpacket : out std_logic;                                        -- startofpacket
			src2_endofpacket   : out std_logic;                                        -- endofpacket
			src3_ready         : in  std_logic                     := 'X';             -- ready
			src3_valid         : out std_logic;                                        -- valid
			src3_data          : out std_logic_vector(93 downto 0);                    -- data
			src3_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src3_startofpacket : out std_logic;                                        -- startofpacket
			src3_endofpacket   : out std_logic;                                        -- endofpacket
			src4_ready         : in  std_logic                     := 'X';             -- ready
			src4_valid         : out std_logic;                                        -- valid
			src4_data          : out std_logic_vector(93 downto 0);                    -- data
			src4_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src4_startofpacket : out std_logic;                                        -- startofpacket
			src4_endofpacket   : out std_logic;                                        -- endofpacket
			src5_ready         : in  std_logic                     := 'X';             -- ready
			src5_valid         : out std_logic;                                        -- valid
			src5_data          : out std_logic_vector(93 downto 0);                    -- data
			src5_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src5_startofpacket : out std_logic;                                        -- startofpacket
			src5_endofpacket   : out std_logic;                                        -- endofpacket
			src6_ready         : in  std_logic                     := 'X';             -- ready
			src6_valid         : out std_logic;                                        -- valid
			src6_data          : out std_logic_vector(93 downto 0);                    -- data
			src6_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src6_startofpacket : out std_logic;                                        -- startofpacket
			src6_endofpacket   : out std_logic;                                        -- endofpacket
			src7_ready         : in  std_logic                     := 'X';             -- ready
			src7_valid         : out std_logic;                                        -- valid
			src7_data          : out std_logic_vector(93 downto 0);                    -- data
			src7_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src7_startofpacket : out std_logic;                                        -- startofpacket
			src7_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component sopc_system_cmd_xbar_demux_007;

	component sopc_system_cmd_xbar_mux_005 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(93 downto 0);                    -- data
			src_channel         : out std_logic_vector(7 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component sopc_system_cmd_xbar_mux_005;

	component sopc_system_rsp_xbar_demux_005 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(93 downto 0);                    -- data
			src0_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(93 downto 0);                    -- data
			src1_channel       : out std_logic_vector(7 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component sopc_system_rsp_xbar_demux_005;

	component sopc_system_rsp_xbar_mux_007 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(93 downto 0);                    -- data
			src_channel         : out std_logic_vector(7 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                        -- ready
			sink2_valid         : in  std_logic                     := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                        -- ready
			sink3_valid         : in  std_logic                     := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink4_ready         : out std_logic;                                        -- ready
			sink4_valid         : in  std_logic                     := 'X';             -- valid
			sink4_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink4_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink4_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink4_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink5_ready         : out std_logic;                                        -- ready
			sink5_valid         : in  std_logic                     := 'X';             -- valid
			sink5_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink5_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink5_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink5_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink6_ready         : out std_logic;                                        -- ready
			sink6_valid         : in  std_logic                     := 'X';             -- valid
			sink6_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink6_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink6_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink6_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink7_ready         : out std_logic;                                        -- ready
			sink7_valid         : in  std_logic                     := 'X';             -- valid
			sink7_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			sink7_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			sink7_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink7_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component sopc_system_rsp_xbar_mux_007;

	component sopc_system_cmd_xbar_demux_008 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- data
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(94 downto 0);                    -- data
			src0_channel       : out std_logic_vector(1 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(94 downto 0);                    -- data
			src1_channel       : out std_logic_vector(1 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component sopc_system_cmd_xbar_demux_008;

	component sopc_system_rsp_xbar_demux_013 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(94 downto 0);                    -- data
			src0_channel       : out std_logic_vector(1 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component sopc_system_rsp_xbar_demux_013;

	component sopc_system_rsp_xbar_mux_008 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(94 downto 0);                    -- data
			src_channel         : out std_logic_vector(1 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component sopc_system_rsp_xbar_mux_008;

	component sopc_system_cmd_xbar_demux_009 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(98 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(98 downto 0);                    -- data
			src0_channel       : out std_logic_vector(1 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component sopc_system_cmd_xbar_demux_009;

	component sopc_system_cmd_xbar_mux_015 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(98 downto 0);                    -- data
			src_channel         : out std_logic_vector(1 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(98 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(98 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component sopc_system_cmd_xbar_mux_015;

	component sopc_system_rsp_xbar_demux_015 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(98 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(98 downto 0);                    -- data
			src0_channel       : out std_logic_vector(1 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(98 downto 0);                    -- data
			src1_channel       : out std_logic_vector(1 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component sopc_system_rsp_xbar_demux_015;

	component sopc_system_cmd_xbar_demux_011 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(96 downto 0);                    -- data
			src0_channel       : out std_logic_vector(1 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component sopc_system_cmd_xbar_demux_011;

	component sopc_system_cmd_xbar_mux_016 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(96 downto 0);                    -- data
			src_channel         : out std_logic_vector(1 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component sopc_system_cmd_xbar_mux_016;

	component sopc_system_rsp_xbar_demux_016 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(96 downto 0);                    -- data
			src0_channel       : out std_logic_vector(1 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(96 downto 0);                    -- data
			src1_channel       : out std_logic_vector(1 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component sopc_system_rsp_xbar_demux_016;

	component sopc_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component sopc_system_irq_mapper;

	component altera_irq_clock_crosser is
		generic (
			IRQ_WIDTH : integer := 1
		);
		port (
			receiver_clk   : in  std_logic                    := 'X';             -- clk
			sender_clk     : in  std_logic                    := 'X';             -- clk
			receiver_reset : in  std_logic                    := 'X';             -- reset
			sender_reset   : in  std_logic                    := 'X';             -- reset
			receiver_irq   : in  std_logic_vector(0 downto 0) := (others => 'X'); -- irq
			sender_irq     : out std_logic_vector(0 downto 0)                     -- irq
		);
	end component altera_irq_clock_crosser;

	component sopc_system_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_ready          : out std_logic;                                        -- ready
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_empty          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			in_0_error          : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- error
			out_0_ready         : in  std_logic                     := 'X';             -- ready
			out_0_valid         : out std_logic;                                        -- valid
			out_0_data          : out std_logic_vector(31 downto 0);                    -- data
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic;                                        -- endofpacket
			out_0_empty         : out std_logic_vector(1 downto 0);                     -- empty
			out_0_error         : out std_logic_vector(5 downto 0)                      -- error
		);
	end component sopc_system_avalon_st_adapter;

	component sopc_system_limiter is
		generic (
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_TRANS_POSTED          : integer := 0;
			PKT_TRANS_WRITE           : integer := 0;
			MAX_OUTSTANDING_RESPONSES : integer := 0;
			PIPELINED                 : integer := 0;
			ST_DATA_W                 : integer := 72;
			ST_CHANNEL_W              : integer := 1;
			VALID_WIDTH               : integer := 1;
			ENFORCE_ORDER             : integer := 1;
			PREVENT_HAZARDS           : integer := 0;
			PKT_BYTE_CNT_H            : integer := 0;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 0;
			PKT_BYTEEN_L              : integer := 0
		);
		port (
			clk                    : in  std_logic                     := 'X';             -- clk
			reset                  : in  std_logic                     := 'X';             -- reset
			cmd_sink_ready         : out std_logic;                                        -- ready
			cmd_sink_valid         : in  std_logic                     := 'X';             -- valid
			cmd_sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			cmd_sink_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			cmd_sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			cmd_sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			cmd_src_ready          : in  std_logic                     := 'X';             -- ready
			cmd_src_data           : out std_logic_vector(99 downto 0);                    -- data
			cmd_src_channel        : out std_logic_vector(3 downto 0);                     -- channel
			cmd_src_startofpacket  : out std_logic;                                        -- startofpacket
			cmd_src_endofpacket    : out std_logic;                                        -- endofpacket
			rsp_sink_ready         : out std_logic;                                        -- ready
			rsp_sink_valid         : in  std_logic                     := 'X';             -- valid
			rsp_sink_channel       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			rsp_sink_data          : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			rsp_sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			rsp_sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			rsp_src_ready          : in  std_logic                     := 'X';             -- ready
			rsp_src_valid          : out std_logic;                                        -- valid
			rsp_src_data           : out std_logic_vector(99 downto 0);                    -- data
			rsp_src_channel        : out std_logic_vector(3 downto 0);                     -- channel
			rsp_src_startofpacket  : out std_logic;                                        -- startofpacket
			rsp_src_endofpacket    : out std_logic;                                        -- endofpacket
			cmd_src_valid          : out std_logic_vector(3 downto 0)                      -- data
		);
	end component sopc_system_limiter;

	component sopc_system_limiter_002 is
		generic (
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_TRANS_POSTED          : integer := 0;
			PKT_TRANS_WRITE           : integer := 0;
			MAX_OUTSTANDING_RESPONSES : integer := 0;
			PIPELINED                 : integer := 0;
			ST_DATA_W                 : integer := 72;
			ST_CHANNEL_W              : integer := 1;
			VALID_WIDTH               : integer := 1;
			ENFORCE_ORDER             : integer := 1;
			PREVENT_HAZARDS           : integer := 0;
			PKT_BYTE_CNT_H            : integer := 0;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 0;
			PKT_BYTEEN_L              : integer := 0
		);
		port (
			clk                    : in  std_logic                     := 'X';             -- clk
			reset                  : in  std_logic                     := 'X';             -- reset
			cmd_sink_ready         : out std_logic;                                        -- ready
			cmd_sink_valid         : in  std_logic                     := 'X';             -- valid
			cmd_sink_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			cmd_sink_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			cmd_sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			cmd_sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			cmd_src_ready          : in  std_logic                     := 'X';             -- ready
			cmd_src_data           : out std_logic_vector(93 downto 0);                    -- data
			cmd_src_channel        : out std_logic_vector(7 downto 0);                     -- channel
			cmd_src_startofpacket  : out std_logic;                                        -- startofpacket
			cmd_src_endofpacket    : out std_logic;                                        -- endofpacket
			rsp_sink_ready         : out std_logic;                                        -- ready
			rsp_sink_valid         : in  std_logic                     := 'X';             -- valid
			rsp_sink_channel       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			rsp_sink_data          : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			rsp_sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			rsp_sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			rsp_src_ready          : in  std_logic                     := 'X';             -- ready
			rsp_src_valid          : out std_logic;                                        -- valid
			rsp_src_data           : out std_logic_vector(93 downto 0);                    -- data
			rsp_src_channel        : out std_logic_vector(7 downto 0);                     -- channel
			rsp_src_startofpacket  : out std_logic;                                        -- startofpacket
			rsp_src_endofpacket    : out std_logic;                                        -- endofpacket
			cmd_src_valid          : out std_logic_vector(7 downto 0)                      -- data
		);
	end component sopc_system_limiter_002;

	component sopc_system_limiter_003 is
		generic (
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_TRANS_POSTED          : integer := 0;
			PKT_TRANS_WRITE           : integer := 0;
			MAX_OUTSTANDING_RESPONSES : integer := 0;
			PIPELINED                 : integer := 0;
			ST_DATA_W                 : integer := 72;
			ST_CHANNEL_W              : integer := 1;
			VALID_WIDTH               : integer := 1;
			ENFORCE_ORDER             : integer := 1;
			PREVENT_HAZARDS           : integer := 0;
			PKT_BYTE_CNT_H            : integer := 0;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 0;
			PKT_BYTEEN_L              : integer := 0
		);
		port (
			clk                    : in  std_logic                     := 'X';             -- clk
			reset                  : in  std_logic                     := 'X';             -- reset
			cmd_sink_ready         : out std_logic;                                        -- ready
			cmd_sink_valid         : in  std_logic                     := 'X';             -- valid
			cmd_sink_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			cmd_sink_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			cmd_sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			cmd_sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			cmd_src_ready          : in  std_logic                     := 'X';             -- ready
			cmd_src_data           : out std_logic_vector(94 downto 0);                    -- data
			cmd_src_channel        : out std_logic_vector(1 downto 0);                     -- channel
			cmd_src_startofpacket  : out std_logic;                                        -- startofpacket
			cmd_src_endofpacket    : out std_logic;                                        -- endofpacket
			rsp_sink_ready         : out std_logic;                                        -- ready
			rsp_sink_valid         : in  std_logic                     := 'X';             -- valid
			rsp_sink_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			rsp_sink_data          : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			rsp_sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			rsp_sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			rsp_src_ready          : in  std_logic                     := 'X';             -- ready
			rsp_src_valid          : out std_logic;                                        -- valid
			rsp_src_data           : out std_logic_vector(94 downto 0);                    -- data
			rsp_src_channel        : out std_logic_vector(1 downto 0);                     -- channel
			rsp_src_startofpacket  : out std_logic;                                        -- startofpacket
			rsp_src_endofpacket    : out std_logic;                                        -- endofpacket
			cmd_src_valid          : out std_logic_vector(1 downto 0)                      -- data
		);
	end component sopc_system_limiter_003;

	component sopc_system_width_adapter is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			in_valid             : in  std_logic                     := 'X';             -- valid
			in_channel           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                     := 'X';             -- endofpacket
			in_ready             : out std_logic;                                        -- ready
			in_data              : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                        -- endofpacket
			out_data             : out std_logic_vector(76 downto 0);                    -- data
			out_channel          : out std_logic_vector(1 downto 0);                     -- channel
			out_valid            : out std_logic;                                        -- valid
			out_ready            : in  std_logic                     := 'X';             -- ready
			out_startofpacket    : out std_logic;                                        -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- data
		);
	end component sopc_system_width_adapter;

	component sopc_system_width_adapter_001 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			in_valid             : in  std_logic                     := 'X';             -- valid
			in_channel           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                     := 'X';             -- endofpacket
			in_ready             : out std_logic;                                        -- ready
			in_data              : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                        -- endofpacket
			out_data             : out std_logic_vector(94 downto 0);                    -- data
			out_channel          : out std_logic_vector(1 downto 0);                     -- channel
			out_valid            : out std_logic;                                        -- valid
			out_ready            : in  std_logic                     := 'X';             -- ready
			out_startofpacket    : out std_logic;                                        -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)  := (others => 'X')  -- data
		);
	end component sopc_system_width_adapter_001;

	component sopc_system_width_adapter_004 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(96 downto 0)  := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(132 downto 0);                    -- data
			out_channel          : out std_logic_vector(1 downto 0);                      -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component sopc_system_width_adapter_004;

	component sopc_system_width_adapter_005 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(132 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(96 downto 0);                     -- data
			out_channel          : out std_logic_vector(1 downto 0);                      -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component sopc_system_width_adapter_005;

	component sopc_system_rst_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component sopc_system_rst_controller;

	component sopc_system_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component sopc_system_rst_controller_002;

	component sopc_system_rst_controller_003 is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component sopc_system_rst_controller_003;

	component sopc_system_rst_controller_004 is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component sopc_system_rst_controller_004;

	component sopc_system_tse_dma_to_sdram_ccb is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			ADDRESS_WIDTH       : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                     := 'X';             -- clk
			m0_reset         : in  std_logic                     := 'X';             -- reset
			s0_clk           : in  std_logic                     := 'X';             -- clk
			s0_reset         : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(26 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component sopc_system_tse_dma_to_sdram_ccb;

	component sopc_system_cpu_to_peripherals_ccb is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			ADDRESS_WIDTH       : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                     := 'X';             -- clk
			m0_reset         : in  std_logic                     := 'X';             -- reset
			s0_clk           : in  std_logic                     := 'X';             -- clk
			s0_reset         : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(22 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(22 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component sopc_system_cpu_to_peripherals_ccb;

	component sopc_system_cpu_to_flash_ccb is
		generic (
			DATA_WIDTH          : integer := 32;
			SYMBOL_WIDTH        : integer := 8;
			ADDRESS_WIDTH       : integer := 10;
			BURSTCOUNT_WIDTH    : integer := 1;
			COMMAND_FIFO_DEPTH  : integer := 4;
			RESPONSE_FIFO_DEPTH : integer := 4;
			MASTER_SYNC_DEPTH   : integer := 2;
			SLAVE_SYNC_DEPTH    : integer := 2
		);
		port (
			m0_clk           : in  std_logic                     := 'X';             -- clk
			m0_reset         : in  std_logic                     := 'X';             -- reset
			s0_clk           : in  std_logic                     := 'X';             -- clk
			s0_reset         : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(27 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component sopc_system_cpu_to_flash_ccb;

	component sopc_system_linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(100 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- address
			csr_read          : in  std_logic                      := 'X';             -- read
			csr_write         : in  std_logic                      := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                         -- data
			almost_empty_data : out std_logic;                                         -- data
			in_empty          : in  std_logic                      := 'X';             -- empty
			out_empty         : out std_logic;                                         -- empty
			in_error          : in  std_logic                      := 'X';             -- error
			out_error         : out std_logic;                                         -- error
			in_channel        : in  std_logic                      := 'X';             -- channel
			out_channel       : out std_logic                                          -- channel
		);
	end component sopc_system_linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component sopc_system_dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(101 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- address
			csr_read          : in  std_logic                      := 'X';             -- read
			csr_write         : in  std_logic                      := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                         -- data
			almost_empty_data : out std_logic;                                         -- data
			in_empty          : in  std_logic                      := 'X';             -- empty
			out_empty         : out std_logic;                                         -- empty
			in_error          : in  std_logic                      := 'X';             -- error
			out_error         : out std_logic;                                         -- error
			in_channel        : in  std_logic                      := 'X';             -- channel
			out_channel       : out std_logic                                          -- channel
		);
	end component sopc_system_dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(94 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component sopc_system_cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(77 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(77 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component sopc_system_cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component sopc_system_cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(17 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component sopc_system_cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component sopc_system_tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(99 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component sopc_system_tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component sopc_system_sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(133 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(133 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- address
			csr_read          : in  std_logic                      := 'X';             -- read
			csr_write         : in  std_logic                      := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                         -- data
			almost_empty_data : out std_logic;                                         -- data
			in_empty          : in  std_logic                      := 'X';             -- empty
			out_empty         : out std_logic;                                         -- empty
			in_error          : in  std_logic                      := 'X';             -- error
			out_error         : out std_logic;                                         -- error
			in_channel        : in  std_logic                      := 'X';             -- channel
			out_channel       : out std_logic                                          -- channel
		);
	end component sopc_system_sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component sopc_system_linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(28 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(99 downto 0);                     -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(99 downto 0)  := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(100 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                         -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                      := 'X'              -- writeresponsevalid
		);
	end component sopc_system_linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent;

	component sopc_system_dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(100 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(101 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                         -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                      := 'X'              -- writeresponsevalid
		);
	end component sopc_system_dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent;

	component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(22 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(93 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(94 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent;

	component sopc_system_cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(27 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(76 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(77 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(77 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(17 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent;

	component sopc_system_tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(31 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(98 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(98 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(99 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent;

	component sopc_system_sdram_0_avl_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(26 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(5 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(7 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(63 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(132 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(132 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(133 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(133 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(65 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(65 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                         -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                      := 'X'              -- writeresponsevalid
		);
	end component sopc_system_sdram_0_avl_translator_avalon_universal_slave_0_agent;

	component sopc_system_linux_cpu_data_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(28 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_linux_cpu_data_master_translator;

	component sopc_system_linux_cpu_instruction_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(28 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_linux_cpu_instruction_master_translator;

	component sopc_system_sgdma_tx_descriptor_write_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_sgdma_tx_descriptor_write_translator;

	component sopc_system_sgdma_rx_descriptor_read_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_sgdma_rx_descriptor_read_translator;

	component sopc_system_dma_to_descriptor_mem_m0_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(22 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_dma_to_descriptor_mem_m0_translator;

	component sopc_system_cpu_to_peripherals_ccb_m0_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(22 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(22 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_cpu_to_peripherals_ccb_m0_translator;

	component sopc_system_cpu_to_flash_ccb_m0_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(27 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_cpu_to_flash_ccb_m0_translator;

	component sopc_system_sgdma_rx_m_write_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(31 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_sgdma_rx_m_write_translator;

	component sopc_system_tse_dma_to_sdram_ccb_m0_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(26 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_tse_dma_to_sdram_ccb_m0_translator;

	component sopc_system_linux_cpu_tightly_coupled_data_master_0_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(28 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_address               : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_clken                 : in  std_logic                     := 'X';             -- clken
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_linux_cpu_tightly_coupled_data_master_0_translator;

	component sopc_system_linux_cpu_tightly_coupled_instruction_master_0_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(28 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_address               : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_clken                 : in  std_logic                     := 'X';             -- clken
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_linux_cpu_tightly_coupled_instruction_master_0_translator;

	component sopc_system_dma_to_descriptor_mem is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			ADDRESS_WIDTH     : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(13 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component sopc_system_dma_to_descriptor_mem;

	component sopc_system_cpu_to_sdram_pb is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			ADDRESS_WIDTH     : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(26 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic                                         -- debugaccess
		);
	end component sopc_system_cpu_to_sdram_pb;

	component sopc_system_linux_cpu_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_linux_cpu_jtag_debug_module_translator;

	component sopc_system_cpu_to_flash_ccb_s0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(27 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_cpu_to_flash_ccb_s0_translator;

	component sopc_system_cpu_to_peripherals_ccb_s0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(22 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_cpu_to_peripherals_ccb_s0_translator;

	component sopc_system_cpu_to_sdram_pb_s0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(26 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_cpu_to_sdram_pb_s0_translator;

	component sopc_system_dma_to_descriptor_mem_s0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(13 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_dma_to_descriptor_mem_s0_translator;

	component sopc_system_descriptor_memory_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(22 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(10 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_descriptor_memory_s1_translator;

	component sopc_system_jtag_uart_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(22 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_jtag_uart_avalon_jtag_slave_translator;

	component sopc_system_tse_mac_control_port_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(22 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(7 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_tse_mac_control_port_translator;

	component sopc_system_sysid_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(22 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_sysid_control_slave_translator;

	component sopc_system_linux_timer_1ms_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(22 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_linux_timer_1ms_s1_translator;

	component sopc_system_gtp_regif_0_s0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(22 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(13 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_gtp_regif_0_s0_translator;

	component sopc_system_sgdma_tx_csr_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(22 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(3 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_sgdma_tx_csr_translator;

	component sopc_system_cfi_flash_ts_controller_fpga_uas_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(26 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_burstcount            : out std_logic_vector(1 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_lock                  : out std_logic;                                        -- lock
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_writebyteenable       : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_cfi_flash_ts_controller_fpga_uas_translator;

	component sopc_system_tse_dma_to_sdram_ccb_s0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(26 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_tse_dma_to_sdram_ccb_s0_translator;

	component sopc_system_sdram_0_avl_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(63 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(23 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(63 downto 0);                    -- writedata
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(2 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(7 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_writebyteenable       : out std_logic_vector(7 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_sdram_0_avl_translator;

	component sopc_system_tlb_miss_ram_1k_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_address               : out std_logic_vector(7 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component sopc_system_tlb_miss_ram_1k_s1_translator;

	component sopc_system_linux_cpu_data_master_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(28 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(99 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(99 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_linux_cpu_data_master_translator_avalon_universal_master_0_agent;

	component sopc_system_sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			av_address              : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- address
			av_write                : in  std_logic                      := 'X';             -- write
			av_read                 : in  std_logic                      := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                     -- readdata
			av_waitrequest          : out std_logic;                                         -- waitrequest
			av_readdatavalid        : out std_logic;                                         -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                      := 'X';             -- debugaccess
			av_lock                 : in  std_logic                      := 'X';             -- lock
			cp_valid                : out std_logic;                                         -- valid
			cp_data                 : out std_logic_vector(100 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_endofpacket          : out std_logic;                                         -- endofpacket
			cp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : in  std_logic                      := 'X';             -- valid
			rp_data                 : in  std_logic_vector(100 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                         -- ready
			av_response             : out std_logic_vector(1 downto 0);                      -- response
			av_writeresponserequest : in  std_logic                      := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                          -- writeresponsevalid
		);
	end component sopc_system_sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent;

	component sopc_system_dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(22 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(93 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(93 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent;

	component sopc_system_cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(94 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(94 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent;

	component sopc_system_sgdma_tx_m_read_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(98 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(98 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_sgdma_tx_m_read_translator_avalon_universal_master_0_agent;

	component sopc_system_tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(96 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(96 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component sopc_system_tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent;

	signal cfi_flash_ts_controller_tcm_chipselect_n_out                                                          : std_logic;                      -- cfi_flash_ts_controller:tcm_chipselect_n_out -> cfi_flash_ts_bridge:tcs_tcm_chipselect_n_out
	signal cfi_flash_ts_controller_tcm_grant                                                                     : std_logic;                      -- cfi_flash_ts_bridge:grant -> cfi_flash_ts_controller:tcm_grant
	signal cfi_flash_ts_controller_tcm_data_outen                                                                : std_logic;                      -- cfi_flash_ts_controller:tcm_data_outen -> cfi_flash_ts_bridge:tcs_tcm_data_outen
	signal cfi_flash_ts_controller_tcm_reset_n_out                                                               : std_logic;                      -- cfi_flash_ts_controller:tcm_reset_n_out -> cfi_flash_ts_bridge:tcs_tcm_reset_n_out
	signal cfi_flash_ts_controller_tcm_outputenable_n_out                                                        : std_logic;                      -- cfi_flash_ts_controller:tcm_outputenable_n_out -> cfi_flash_ts_bridge:tcs_tcm_outputenable_n_out
	signal cfi_flash_ts_controller_tcm_request                                                                   : std_logic;                      -- cfi_flash_ts_controller:tcm_request -> cfi_flash_ts_bridge:request
	signal cfi_flash_ts_controller_tcm_data_out                                                                  : std_logic_vector(15 downto 0);  -- cfi_flash_ts_controller:tcm_data_out -> cfi_flash_ts_bridge:tcs_tcm_data_out
	signal cfi_flash_ts_controller_tcm_write_n_out                                                               : std_logic;                      -- cfi_flash_ts_controller:tcm_write_n_out -> cfi_flash_ts_bridge:tcs_tcm_write_n_out
	signal cfi_flash_ts_controller_tcm_address_out                                                               : std_logic_vector(26 downto 0);  -- cfi_flash_ts_controller:tcm_address_out -> cfi_flash_ts_bridge:tcs_tcm_address_out
	signal cfi_flash_ts_controller_tcm_data_in                                                                   : std_logic_vector(15 downto 0);  -- cfi_flash_ts_bridge:tcs_tcm_data_in -> cfi_flash_ts_controller:tcm_data_in
	signal sgdma_tx_out_endofpacket                                                                              : std_logic;                      -- sgdma_tx:out_endofpacket -> tse_mac:ff_tx_eop
	signal sgdma_tx_out_valid                                                                                    : std_logic;                      -- sgdma_tx:out_valid -> tse_mac:ff_tx_wren
	signal sgdma_tx_out_startofpacket                                                                            : std_logic;                      -- sgdma_tx:out_startofpacket -> tse_mac:ff_tx_sop
	signal sgdma_tx_out_error                                                                                    : std_logic;                      -- sgdma_tx:out_error -> tse_mac:ff_tx_err
	signal sgdma_tx_out_empty                                                                                    : std_logic_vector(1 downto 0);   -- sgdma_tx:out_empty -> tse_mac:ff_tx_mod
	signal sgdma_tx_out_data                                                                                     : std_logic_vector(31 downto 0);  -- sgdma_tx:out_data -> tse_mac:ff_tx_data
	signal sgdma_tx_out_ready                                                                                    : std_logic;                      -- tse_mac:ff_tx_rdy -> sgdma_tx:out_ready
	signal cfi_flash_ts_controller_fpga_tcm_chipselect_n_out                                                     : std_logic;                      -- cfi_flash_ts_controller_fpga:tcm_chipselect_n_out -> cfi_flash_ts_bridge_fpga:tcs_tcm_chipselect_n_out
	signal cfi_flash_ts_controller_fpga_tcm_grant                                                                : std_logic;                      -- cfi_flash_ts_bridge_fpga:grant -> cfi_flash_ts_controller_fpga:tcm_grant
	signal cfi_flash_ts_controller_fpga_tcm_data_outen                                                           : std_logic;                      -- cfi_flash_ts_controller_fpga:tcm_data_outen -> cfi_flash_ts_bridge_fpga:tcs_tcm_data_outen
	signal cfi_flash_ts_controller_fpga_tcm_reset_n_out                                                          : std_logic;                      -- cfi_flash_ts_controller_fpga:tcm_reset_n_out -> cfi_flash_ts_bridge_fpga:tcs_tcm_reset_n_out
	signal cfi_flash_ts_controller_fpga_tcm_outputenable_n_out                                                   : std_logic;                      -- cfi_flash_ts_controller_fpga:tcm_outputenable_n_out -> cfi_flash_ts_bridge_fpga:tcs_tcm_outputenable_n_out
	signal cfi_flash_ts_controller_fpga_tcm_request                                                              : std_logic;                      -- cfi_flash_ts_controller_fpga:tcm_request -> cfi_flash_ts_bridge_fpga:request
	signal cfi_flash_ts_controller_fpga_tcm_data_out                                                             : std_logic_vector(15 downto 0);  -- cfi_flash_ts_controller_fpga:tcm_data_out -> cfi_flash_ts_bridge_fpga:tcs_tcm_data_out
	signal cfi_flash_ts_controller_fpga_tcm_write_n_out                                                          : std_logic;                      -- cfi_flash_ts_controller_fpga:tcm_write_n_out -> cfi_flash_ts_bridge_fpga:tcs_tcm_write_n_out
	signal cfi_flash_ts_controller_fpga_tcm_address_out                                                          : std_logic_vector(26 downto 0);  -- cfi_flash_ts_controller_fpga:tcm_address_out -> cfi_flash_ts_bridge_fpga:tcs_tcm_address_out
	signal cfi_flash_ts_controller_fpga_tcm_data_in                                                              : std_logic_vector(15 downto 0);  -- cfi_flash_ts_bridge_fpga:tcs_tcm_data_in -> cfi_flash_ts_controller_fpga:tcm_data_in
	signal sdram_0_afi_clk_clk                                                                                   : std_logic;                      -- sdram_0:afi_clk -> [addr_router:clk, addr_router_001:clk, addr_router_011:clk, addr_router_012:clk, cmd_xbar_demux:clk, cmd_xbar_demux_001:clk, cmd_xbar_demux_011:clk, cmd_xbar_demux_012:clk, cmd_xbar_mux:clk, cmd_xbar_mux_001:clk, cmd_xbar_mux_003:clk, cmd_xbar_mux_016:clk, cpu_to_flash_ccb:s0_clk, cpu_to_flash_ccb_s0_translator:clk, cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:clk, cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cpu_to_peripherals_ccb:s0_clk, cpu_to_peripherals_ccb_s0_translator:clk, cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:clk, cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cpu_to_sdram_pb:clk, cpu_to_sdram_pb_m0_translator:clk, cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:clk, cpu_to_sdram_pb_s0_translator:clk, cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:clk, cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, id_router_016:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, irq_synchronizer_003:sender_clk, irq_synchronizer_004:sender_clk, limiter:clk, limiter_001:clk, linux_cpu:clk, linux_cpu_data_master_translator:clk, linux_cpu_data_master_translator_avalon_universal_master_0_agent:clk, linux_cpu_instruction_master_translator:clk, linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:clk, linux_cpu_jtag_debug_module_translator:clk, linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:clk, linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, linux_cpu_tightly_coupled_data_master_0_translator:clk, linux_cpu_tightly_coupled_instruction_master_0_translator:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_demux_016:clk, rsp_xbar_mux:clk, rsp_xbar_mux_001:clk, rst_controller_001:clk, rst_controller_004:clk, sdram_0_avl_translator:clk, sdram_0_avl_translator_avalon_universal_slave_0_agent:clk, sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, tlb_miss_ram_1k:clk, tlb_miss_ram_1k:clk2, tlb_miss_ram_1k_s1_translator:clk, tlb_miss_ram_1k_s2_translator:clk, tse_dma_to_sdram_ccb:m0_clk, tse_dma_to_sdram_ccb_m0_translator:clk, tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:clk, width_adapter_004:clk, width_adapter_005:clk]
	signal sdram_0_afi_half_clk_clk                                                                              : std_logic;                      -- sdram_0:afi_half_clk -> [addr_router_002:clk, addr_router_003:clk, addr_router_004:clk, addr_router_005:clk, addr_router_006:clk, addr_router_007:clk, addr_router_008:clk, addr_router_009:clk, addr_router_010:clk, avalon_st_adapter:in_clk_0_clk, burst_adapter:clk, burst_adapter_001:clk, cfi_flash_ts_bridge:clk, cfi_flash_ts_bridge_fpga:clk, cfi_flash_ts_controller:clk_clk, cfi_flash_ts_controller_fpga:clk_clk, cfi_flash_ts_controller_fpga_uas_translator:clk, cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:clk, cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cfi_flash_ts_controller_uas_translator:clk, cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:clk, cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, cmd_xbar_demux_002:clk, cmd_xbar_demux_003:clk, cmd_xbar_demux_004:clk, cmd_xbar_demux_005:clk, cmd_xbar_demux_006:clk, cmd_xbar_demux_007:clk, cmd_xbar_demux_008:clk, cmd_xbar_demux_009:clk, cmd_xbar_demux_010:clk, cmd_xbar_mux_004:clk, cmd_xbar_mux_005:clk, cmd_xbar_mux_015:clk, cpu_to_flash_ccb:m0_clk, cpu_to_flash_ccb_m0_translator:clk, cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:clk, cpu_to_peripherals_ccb:m0_clk, cpu_to_peripherals_ccb_m0_translator:clk, cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:clk, descriptor_memory:clk, descriptor_memory_s1_translator:clk, descriptor_memory_s1_translator_avalon_universal_slave_0_agent:clk, descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, dma_to_descriptor_mem:clk, dma_to_descriptor_mem_m0_translator:clk, dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:clk, dma_to_descriptor_mem_s0_translator:clk, dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:clk, dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, gtp_regif_0:clk, gtp_regif_0_s0_translator:clk, gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:clk, gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router_004:clk, id_router_005:clk, id_router_006:clk, id_router_007:clk, id_router_008:clk, id_router_009:clk, id_router_010:clk, id_router_011:clk, id_router_012:clk, id_router_013:clk, id_router_014:clk, id_router_015:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_002:receiver_clk, irq_synchronizer_003:receiver_clk, irq_synchronizer_004:receiver_clk, jtag_uart:clk, jtag_uart_avalon_jtag_slave_translator:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:clk, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, limiter_002:clk, limiter_003:clk, linux_timer_1ms:clk, linux_timer_1ms_s1_translator:clk, linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:clk, linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux_004:clk, rsp_xbar_demux_005:clk, rsp_xbar_demux_006:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rsp_xbar_demux_009:clk, rsp_xbar_demux_010:clk, rsp_xbar_demux_011:clk, rsp_xbar_demux_012:clk, rsp_xbar_demux_013:clk, rsp_xbar_demux_014:clk, rsp_xbar_demux_015:clk, rsp_xbar_mux_007:clk, rsp_xbar_mux_008:clk, rst_controller:clk, rst_controller_003:clk, sgdma_rx:clk, sgdma_rx_csr_translator:clk, sgdma_rx_csr_translator_avalon_universal_slave_0_agent:clk, sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sgdma_rx_descriptor_read_translator:clk, sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:clk, sgdma_rx_descriptor_write_translator:clk, sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:clk, sgdma_rx_m_write_translator:clk, sgdma_rx_m_write_translator_avalon_universal_master_0_agent:clk, sgdma_tx:clk, sgdma_tx_csr_translator:clk, sgdma_tx_csr_translator_avalon_universal_slave_0_agent:clk, sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, sgdma_tx_descriptor_read_translator:clk, sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:clk, sgdma_tx_descriptor_write_translator:clk, sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:clk, sgdma_tx_m_read_translator:clk, sgdma_tx_m_read_translator_avalon_universal_master_0_agent:clk, sysid:clock, sysid_control_slave_translator:clk, sysid_control_slave_translator_avalon_universal_slave_0_agent:clk, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, tse_dma_to_sdram_ccb:s0_clk, tse_dma_to_sdram_ccb_s0_translator:clk, tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:clk, tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, tse_mac:clk, tse_mac:ff_rx_clk, tse_mac:ff_tx_clk, tse_mac_control_port_translator:clk, tse_mac_control_port_translator_avalon_universal_slave_0_agent:clk, tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk]
	signal linux_cpu_data_master_waitrequest                                                                     : std_logic;                      -- linux_cpu_data_master_translator:av_waitrequest -> linux_cpu:d_waitrequest
	signal linux_cpu_data_master_writedata                                                                       : std_logic_vector(31 downto 0);  -- linux_cpu:d_writedata -> linux_cpu_data_master_translator:av_writedata
	signal linux_cpu_data_master_address                                                                         : std_logic_vector(28 downto 0);  -- linux_cpu:d_address -> linux_cpu_data_master_translator:av_address
	signal linux_cpu_data_master_write                                                                           : std_logic;                      -- linux_cpu:d_write -> linux_cpu_data_master_translator:av_write
	signal linux_cpu_data_master_read                                                                            : std_logic;                      -- linux_cpu:d_read -> linux_cpu_data_master_translator:av_read
	signal linux_cpu_data_master_readdata                                                                        : std_logic_vector(31 downto 0);  -- linux_cpu_data_master_translator:av_readdata -> linux_cpu:d_readdata
	signal linux_cpu_data_master_debugaccess                                                                     : std_logic;                      -- linux_cpu:jtag_debug_module_debugaccess_to_roms -> linux_cpu_data_master_translator:av_debugaccess
	signal linux_cpu_data_master_readdatavalid                                                                   : std_logic;                      -- linux_cpu_data_master_translator:av_readdatavalid -> linux_cpu:d_readdatavalid
	signal linux_cpu_data_master_byteenable                                                                      : std_logic_vector(3 downto 0);   -- linux_cpu:d_byteenable -> linux_cpu_data_master_translator:av_byteenable
	signal linux_cpu_instruction_master_waitrequest                                                              : std_logic;                      -- linux_cpu_instruction_master_translator:av_waitrequest -> linux_cpu:i_waitrequest
	signal linux_cpu_instruction_master_address                                                                  : std_logic_vector(28 downto 0);  -- linux_cpu:i_address -> linux_cpu_instruction_master_translator:av_address
	signal linux_cpu_instruction_master_read                                                                     : std_logic;                      -- linux_cpu:i_read -> linux_cpu_instruction_master_translator:av_read
	signal linux_cpu_instruction_master_readdata                                                                 : std_logic_vector(31 downto 0);  -- linux_cpu_instruction_master_translator:av_readdata -> linux_cpu:i_readdata
	signal linux_cpu_instruction_master_readdatavalid                                                            : std_logic;                      -- linux_cpu_instruction_master_translator:av_readdatavalid -> linux_cpu:i_readdatavalid
	signal linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest                                : std_logic;                      -- linux_cpu:jtag_debug_module_waitrequest -> linux_cpu_jtag_debug_module_translator:av_waitrequest
	signal linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata                                  : std_logic_vector(31 downto 0);  -- linux_cpu_jtag_debug_module_translator:av_writedata -> linux_cpu:jtag_debug_module_writedata
	signal linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_address                                    : std_logic_vector(8 downto 0);   -- linux_cpu_jtag_debug_module_translator:av_address -> linux_cpu:jtag_debug_module_address
	signal linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_write                                      : std_logic;                      -- linux_cpu_jtag_debug_module_translator:av_write -> linux_cpu:jtag_debug_module_write
	signal linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_read                                       : std_logic;                      -- linux_cpu_jtag_debug_module_translator:av_read -> linux_cpu:jtag_debug_module_read
	signal linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata                                   : std_logic_vector(31 downto 0);  -- linux_cpu:jtag_debug_module_readdata -> linux_cpu_jtag_debug_module_translator:av_readdata
	signal linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                                : std_logic;                      -- linux_cpu_jtag_debug_module_translator:av_debugaccess -> linux_cpu:jtag_debug_module_debugaccess
	signal linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                                 : std_logic_vector(3 downto 0);   -- linux_cpu_jtag_debug_module_translator:av_byteenable -> linux_cpu:jtag_debug_module_byteenable
	signal cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_waitrequest                                        : std_logic;                      -- cpu_to_flash_ccb:s0_waitrequest -> cpu_to_flash_ccb_s0_translator:av_waitrequest
	signal cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_burstcount                                         : std_logic_vector(0 downto 0);   -- cpu_to_flash_ccb_s0_translator:av_burstcount -> cpu_to_flash_ccb:s0_burstcount
	signal cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_writedata                                          : std_logic_vector(31 downto 0);  -- cpu_to_flash_ccb_s0_translator:av_writedata -> cpu_to_flash_ccb:s0_writedata
	signal cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_address                                            : std_logic_vector(27 downto 0);  -- cpu_to_flash_ccb_s0_translator:av_address -> cpu_to_flash_ccb:s0_address
	signal cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_write                                              : std_logic;                      -- cpu_to_flash_ccb_s0_translator:av_write -> cpu_to_flash_ccb:s0_write
	signal cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_read                                               : std_logic;                      -- cpu_to_flash_ccb_s0_translator:av_read -> cpu_to_flash_ccb:s0_read
	signal cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_readdata                                           : std_logic_vector(31 downto 0);  -- cpu_to_flash_ccb:s0_readdata -> cpu_to_flash_ccb_s0_translator:av_readdata
	signal cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_debugaccess                                        : std_logic;                      -- cpu_to_flash_ccb_s0_translator:av_debugaccess -> cpu_to_flash_ccb:s0_debugaccess
	signal cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_readdatavalid                                      : std_logic;                      -- cpu_to_flash_ccb:s0_readdatavalid -> cpu_to_flash_ccb_s0_translator:av_readdatavalid
	signal cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_byteenable                                         : std_logic_vector(3 downto 0);   -- cpu_to_flash_ccb_s0_translator:av_byteenable -> cpu_to_flash_ccb:s0_byteenable
	signal cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_waitrequest                                  : std_logic;                      -- cpu_to_peripherals_ccb:s0_waitrequest -> cpu_to_peripherals_ccb_s0_translator:av_waitrequest
	signal cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_burstcount                                   : std_logic_vector(0 downto 0);   -- cpu_to_peripherals_ccb_s0_translator:av_burstcount -> cpu_to_peripherals_ccb:s0_burstcount
	signal cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_writedata                                    : std_logic_vector(31 downto 0);  -- cpu_to_peripherals_ccb_s0_translator:av_writedata -> cpu_to_peripherals_ccb:s0_writedata
	signal cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_address                                      : std_logic_vector(22 downto 0);  -- cpu_to_peripherals_ccb_s0_translator:av_address -> cpu_to_peripherals_ccb:s0_address
	signal cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_write                                        : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator:av_write -> cpu_to_peripherals_ccb:s0_write
	signal cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_read                                         : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator:av_read -> cpu_to_peripherals_ccb:s0_read
	signal cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_readdata                                     : std_logic_vector(31 downto 0);  -- cpu_to_peripherals_ccb:s0_readdata -> cpu_to_peripherals_ccb_s0_translator:av_readdata
	signal cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_debugaccess                                  : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator:av_debugaccess -> cpu_to_peripherals_ccb:s0_debugaccess
	signal cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_readdatavalid                                : std_logic;                      -- cpu_to_peripherals_ccb:s0_readdatavalid -> cpu_to_peripherals_ccb_s0_translator:av_readdatavalid
	signal cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_byteenable                                   : std_logic_vector(3 downto 0);   -- cpu_to_peripherals_ccb_s0_translator:av_byteenable -> cpu_to_peripherals_ccb:s0_byteenable
	signal cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_waitrequest                                         : std_logic;                      -- cpu_to_sdram_pb:s0_waitrequest -> cpu_to_sdram_pb_s0_translator:av_waitrequest
	signal cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_burstcount                                          : std_logic_vector(0 downto 0);   -- cpu_to_sdram_pb_s0_translator:av_burstcount -> cpu_to_sdram_pb:s0_burstcount
	signal cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_writedata                                           : std_logic_vector(31 downto 0);  -- cpu_to_sdram_pb_s0_translator:av_writedata -> cpu_to_sdram_pb:s0_writedata
	signal cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_address                                             : std_logic_vector(26 downto 0);  -- cpu_to_sdram_pb_s0_translator:av_address -> cpu_to_sdram_pb:s0_address
	signal cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_write                                               : std_logic;                      -- cpu_to_sdram_pb_s0_translator:av_write -> cpu_to_sdram_pb:s0_write
	signal cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_read                                                : std_logic;                      -- cpu_to_sdram_pb_s0_translator:av_read -> cpu_to_sdram_pb:s0_read
	signal cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_readdata                                            : std_logic_vector(31 downto 0);  -- cpu_to_sdram_pb:s0_readdata -> cpu_to_sdram_pb_s0_translator:av_readdata
	signal cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_debugaccess                                         : std_logic;                      -- cpu_to_sdram_pb_s0_translator:av_debugaccess -> cpu_to_sdram_pb:s0_debugaccess
	signal cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_readdatavalid                                       : std_logic;                      -- cpu_to_sdram_pb:s0_readdatavalid -> cpu_to_sdram_pb_s0_translator:av_readdatavalid
	signal cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_byteenable                                          : std_logic_vector(3 downto 0);   -- cpu_to_sdram_pb_s0_translator:av_byteenable -> cpu_to_sdram_pb:s0_byteenable
	signal sgdma_tx_descriptor_write_waitrequest                                                                 : std_logic;                      -- sgdma_tx_descriptor_write_translator:av_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	signal sgdma_tx_descriptor_write_writedata                                                                   : std_logic_vector(31 downto 0);  -- sgdma_tx:descriptor_write_writedata -> sgdma_tx_descriptor_write_translator:av_writedata
	signal sgdma_tx_descriptor_write_address                                                                     : std_logic_vector(31 downto 0);  -- sgdma_tx:descriptor_write_address -> sgdma_tx_descriptor_write_translator:av_address
	signal sgdma_tx_descriptor_write_write                                                                       : std_logic;                      -- sgdma_tx:descriptor_write_write -> sgdma_tx_descriptor_write_translator:av_write
	signal sgdma_rx_descriptor_write_waitrequest                                                                 : std_logic;                      -- sgdma_rx_descriptor_write_translator:av_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	signal sgdma_rx_descriptor_write_writedata                                                                   : std_logic_vector(31 downto 0);  -- sgdma_rx:descriptor_write_writedata -> sgdma_rx_descriptor_write_translator:av_writedata
	signal sgdma_rx_descriptor_write_address                                                                     : std_logic_vector(31 downto 0);  -- sgdma_rx:descriptor_write_address -> sgdma_rx_descriptor_write_translator:av_address
	signal sgdma_rx_descriptor_write_write                                                                       : std_logic;                      -- sgdma_rx:descriptor_write_write -> sgdma_rx_descriptor_write_translator:av_write
	signal sgdma_rx_descriptor_read_waitrequest                                                                  : std_logic;                      -- sgdma_rx_descriptor_read_translator:av_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	signal sgdma_rx_descriptor_read_address                                                                      : std_logic_vector(31 downto 0);  -- sgdma_rx:descriptor_read_address -> sgdma_rx_descriptor_read_translator:av_address
	signal sgdma_rx_descriptor_read_read                                                                         : std_logic;                      -- sgdma_rx:descriptor_read_read -> sgdma_rx_descriptor_read_translator:av_read
	signal sgdma_rx_descriptor_read_readdata                                                                     : std_logic_vector(31 downto 0);  -- sgdma_rx_descriptor_read_translator:av_readdata -> sgdma_rx:descriptor_read_readdata
	signal sgdma_rx_descriptor_read_readdatavalid                                                                : std_logic;                      -- sgdma_rx_descriptor_read_translator:av_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	signal sgdma_tx_descriptor_read_waitrequest                                                                  : std_logic;                      -- sgdma_tx_descriptor_read_translator:av_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	signal sgdma_tx_descriptor_read_address                                                                      : std_logic_vector(31 downto 0);  -- sgdma_tx:descriptor_read_address -> sgdma_tx_descriptor_read_translator:av_address
	signal sgdma_tx_descriptor_read_read                                                                         : std_logic;                      -- sgdma_tx:descriptor_read_read -> sgdma_tx_descriptor_read_translator:av_read
	signal sgdma_tx_descriptor_read_readdata                                                                     : std_logic_vector(31 downto 0);  -- sgdma_tx_descriptor_read_translator:av_readdata -> sgdma_tx:descriptor_read_readdata
	signal sgdma_tx_descriptor_read_readdatavalid                                                                : std_logic;                      -- sgdma_tx_descriptor_read_translator:av_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	signal dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_waitrequest                                   : std_logic;                      -- dma_to_descriptor_mem:s0_waitrequest -> dma_to_descriptor_mem_s0_translator:av_waitrequest
	signal dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_burstcount                                    : std_logic_vector(0 downto 0);   -- dma_to_descriptor_mem_s0_translator:av_burstcount -> dma_to_descriptor_mem:s0_burstcount
	signal dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_writedata                                     : std_logic_vector(31 downto 0);  -- dma_to_descriptor_mem_s0_translator:av_writedata -> dma_to_descriptor_mem:s0_writedata
	signal dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_address                                       : std_logic_vector(13 downto 0);  -- dma_to_descriptor_mem_s0_translator:av_address -> dma_to_descriptor_mem:s0_address
	signal dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_write                                         : std_logic;                      -- dma_to_descriptor_mem_s0_translator:av_write -> dma_to_descriptor_mem:s0_write
	signal dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_read                                          : std_logic;                      -- dma_to_descriptor_mem_s0_translator:av_read -> dma_to_descriptor_mem:s0_read
	signal dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_readdata                                      : std_logic_vector(31 downto 0);  -- dma_to_descriptor_mem:s0_readdata -> dma_to_descriptor_mem_s0_translator:av_readdata
	signal dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_debugaccess                                   : std_logic;                      -- dma_to_descriptor_mem_s0_translator:av_debugaccess -> dma_to_descriptor_mem:s0_debugaccess
	signal dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_readdatavalid                                 : std_logic;                      -- dma_to_descriptor_mem:s0_readdatavalid -> dma_to_descriptor_mem_s0_translator:av_readdatavalid
	signal dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_byteenable                                    : std_logic_vector(3 downto 0);   -- dma_to_descriptor_mem_s0_translator:av_byteenable -> dma_to_descriptor_mem:s0_byteenable
	signal dma_to_descriptor_mem_m0_burstcount                                                                   : std_logic_vector(0 downto 0);   -- dma_to_descriptor_mem:m0_burstcount -> dma_to_descriptor_mem_m0_translator:av_burstcount
	signal dma_to_descriptor_mem_m0_waitrequest                                                                  : std_logic;                      -- dma_to_descriptor_mem_m0_translator:av_waitrequest -> dma_to_descriptor_mem:m0_waitrequest
	signal dma_to_descriptor_mem_m0_address                                                                      : std_logic_vector(13 downto 0);  -- dma_to_descriptor_mem:m0_address -> dma_to_descriptor_mem_m0_translator:av_address
	signal dma_to_descriptor_mem_m0_writedata                                                                    : std_logic_vector(31 downto 0);  -- dma_to_descriptor_mem:m0_writedata -> dma_to_descriptor_mem_m0_translator:av_writedata
	signal dma_to_descriptor_mem_m0_write                                                                        : std_logic;                      -- dma_to_descriptor_mem:m0_write -> dma_to_descriptor_mem_m0_translator:av_write
	signal dma_to_descriptor_mem_m0_read                                                                         : std_logic;                      -- dma_to_descriptor_mem:m0_read -> dma_to_descriptor_mem_m0_translator:av_read
	signal dma_to_descriptor_mem_m0_readdata                                                                     : std_logic_vector(31 downto 0);  -- dma_to_descriptor_mem_m0_translator:av_readdata -> dma_to_descriptor_mem:m0_readdata
	signal dma_to_descriptor_mem_m0_debugaccess                                                                  : std_logic;                      -- dma_to_descriptor_mem:m0_debugaccess -> dma_to_descriptor_mem_m0_translator:av_debugaccess
	signal dma_to_descriptor_mem_m0_byteenable                                                                   : std_logic_vector(3 downto 0);   -- dma_to_descriptor_mem:m0_byteenable -> dma_to_descriptor_mem_m0_translator:av_byteenable
	signal dma_to_descriptor_mem_m0_readdatavalid                                                                : std_logic;                      -- dma_to_descriptor_mem_m0_translator:av_readdatavalid -> dma_to_descriptor_mem:m0_readdatavalid
	signal cpu_to_peripherals_ccb_m0_burstcount                                                                  : std_logic_vector(0 downto 0);   -- cpu_to_peripherals_ccb:m0_burstcount -> cpu_to_peripherals_ccb_m0_translator:av_burstcount
	signal cpu_to_peripherals_ccb_m0_waitrequest                                                                 : std_logic;                      -- cpu_to_peripherals_ccb_m0_translator:av_waitrequest -> cpu_to_peripherals_ccb:m0_waitrequest
	signal cpu_to_peripherals_ccb_m0_address                                                                     : std_logic_vector(22 downto 0);  -- cpu_to_peripherals_ccb:m0_address -> cpu_to_peripherals_ccb_m0_translator:av_address
	signal cpu_to_peripherals_ccb_m0_writedata                                                                   : std_logic_vector(31 downto 0);  -- cpu_to_peripherals_ccb:m0_writedata -> cpu_to_peripherals_ccb_m0_translator:av_writedata
	signal cpu_to_peripherals_ccb_m0_write                                                                       : std_logic;                      -- cpu_to_peripherals_ccb:m0_write -> cpu_to_peripherals_ccb_m0_translator:av_write
	signal cpu_to_peripherals_ccb_m0_read                                                                        : std_logic;                      -- cpu_to_peripherals_ccb:m0_read -> cpu_to_peripherals_ccb_m0_translator:av_read
	signal cpu_to_peripherals_ccb_m0_readdata                                                                    : std_logic_vector(31 downto 0);  -- cpu_to_peripherals_ccb_m0_translator:av_readdata -> cpu_to_peripherals_ccb:m0_readdata
	signal cpu_to_peripherals_ccb_m0_debugaccess                                                                 : std_logic;                      -- cpu_to_peripherals_ccb:m0_debugaccess -> cpu_to_peripherals_ccb_m0_translator:av_debugaccess
	signal cpu_to_peripherals_ccb_m0_byteenable                                                                  : std_logic_vector(3 downto 0);   -- cpu_to_peripherals_ccb:m0_byteenable -> cpu_to_peripherals_ccb_m0_translator:av_byteenable
	signal cpu_to_peripherals_ccb_m0_readdatavalid                                                               : std_logic;                      -- cpu_to_peripherals_ccb_m0_translator:av_readdatavalid -> cpu_to_peripherals_ccb:m0_readdatavalid
	signal descriptor_memory_s1_translator_avalon_anti_slave_0_writedata                                         : std_logic_vector(31 downto 0);  -- descriptor_memory_s1_translator:av_writedata -> descriptor_memory:writedata
	signal descriptor_memory_s1_translator_avalon_anti_slave_0_address                                           : std_logic_vector(10 downto 0);  -- descriptor_memory_s1_translator:av_address -> descriptor_memory:address
	signal descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect                                        : std_logic;                      -- descriptor_memory_s1_translator:av_chipselect -> descriptor_memory:chipselect
	signal descriptor_memory_s1_translator_avalon_anti_slave_0_clken                                             : std_logic;                      -- descriptor_memory_s1_translator:av_clken -> descriptor_memory:clken
	signal descriptor_memory_s1_translator_avalon_anti_slave_0_write                                             : std_logic;                      -- descriptor_memory_s1_translator:av_write -> descriptor_memory:write
	signal descriptor_memory_s1_translator_avalon_anti_slave_0_readdata                                          : std_logic_vector(31 downto 0);  -- descriptor_memory:readdata -> descriptor_memory_s1_translator:av_readdata
	signal descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable                                        : std_logic_vector(3 downto 0);   -- descriptor_memory_s1_translator:av_byteenable -> descriptor_memory:byteenable
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                                : std_logic;                      -- jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                                  : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                    : std_logic_vector(0 downto 0);   -- jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                                 : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                      : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                       : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                                   : std_logic_vector(31 downto 0);  -- jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	signal tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest                                       : std_logic;                      -- tse_mac:waitrequest -> tse_mac_control_port_translator:av_waitrequest
	signal tse_mac_control_port_translator_avalon_anti_slave_0_writedata                                         : std_logic_vector(31 downto 0);  -- tse_mac_control_port_translator:av_writedata -> tse_mac:writedata
	signal tse_mac_control_port_translator_avalon_anti_slave_0_address                                           : std_logic_vector(7 downto 0);   -- tse_mac_control_port_translator:av_address -> tse_mac:address
	signal tse_mac_control_port_translator_avalon_anti_slave_0_write                                             : std_logic;                      -- tse_mac_control_port_translator:av_write -> tse_mac:write
	signal tse_mac_control_port_translator_avalon_anti_slave_0_read                                              : std_logic;                      -- tse_mac_control_port_translator:av_read -> tse_mac:read
	signal tse_mac_control_port_translator_avalon_anti_slave_0_readdata                                          : std_logic_vector(31 downto 0);  -- tse_mac:readdata -> tse_mac_control_port_translator:av_readdata
	signal sysid_control_slave_translator_avalon_anti_slave_0_address                                            : std_logic_vector(0 downto 0);   -- sysid_control_slave_translator:av_address -> sysid:address
	signal sysid_control_slave_translator_avalon_anti_slave_0_readdata                                           : std_logic_vector(31 downto 0);  -- sysid:readdata -> sysid_control_slave_translator:av_readdata
	signal linux_timer_1ms_s1_translator_avalon_anti_slave_0_writedata                                           : std_logic_vector(15 downto 0);  -- linux_timer_1ms_s1_translator:av_writedata -> linux_timer_1ms:writedata
	signal linux_timer_1ms_s1_translator_avalon_anti_slave_0_address                                             : std_logic_vector(2 downto 0);   -- linux_timer_1ms_s1_translator:av_address -> linux_timer_1ms:address
	signal linux_timer_1ms_s1_translator_avalon_anti_slave_0_chipselect                                          : std_logic;                      -- linux_timer_1ms_s1_translator:av_chipselect -> linux_timer_1ms:chipselect
	signal linux_timer_1ms_s1_translator_avalon_anti_slave_0_write                                               : std_logic;                      -- linux_timer_1ms_s1_translator:av_write -> linux_timer_1ms_s1_translator_avalon_anti_slave_0_write:in
	signal linux_timer_1ms_s1_translator_avalon_anti_slave_0_readdata                                            : std_logic_vector(15 downto 0);  -- linux_timer_1ms:readdata -> linux_timer_1ms_s1_translator:av_readdata
	signal gtp_regif_0_s0_translator_avalon_anti_slave_0_waitrequest                                             : std_logic;                      -- gtp_regif_0:avs_s0_waitrequest -> gtp_regif_0_s0_translator:av_waitrequest
	signal gtp_regif_0_s0_translator_avalon_anti_slave_0_writedata                                               : std_logic_vector(31 downto 0);  -- gtp_regif_0_s0_translator:av_writedata -> gtp_regif_0:avs_s0_writedata
	signal gtp_regif_0_s0_translator_avalon_anti_slave_0_address                                                 : std_logic_vector(13 downto 0);  -- gtp_regif_0_s0_translator:av_address -> gtp_regif_0:avs_s0_address
	signal gtp_regif_0_s0_translator_avalon_anti_slave_0_write                                                   : std_logic;                      -- gtp_regif_0_s0_translator:av_write -> gtp_regif_0:avs_s0_write
	signal gtp_regif_0_s0_translator_avalon_anti_slave_0_read                                                    : std_logic;                      -- gtp_regif_0_s0_translator:av_read -> gtp_regif_0:avs_s0_read
	signal gtp_regif_0_s0_translator_avalon_anti_slave_0_readdata                                                : std_logic_vector(31 downto 0);  -- gtp_regif_0:avs_s0_readdata -> gtp_regif_0_s0_translator:av_readdata
	signal sgdma_tx_csr_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(31 downto 0);  -- sgdma_tx_csr_translator:av_writedata -> sgdma_tx:csr_writedata
	signal sgdma_tx_csr_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(3 downto 0);   -- sgdma_tx_csr_translator:av_address -> sgdma_tx:csr_address
	signal sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect                                                : std_logic;                      -- sgdma_tx_csr_translator:av_chipselect -> sgdma_tx:csr_chipselect
	signal sgdma_tx_csr_translator_avalon_anti_slave_0_write                                                     : std_logic;                      -- sgdma_tx_csr_translator:av_write -> sgdma_tx:csr_write
	signal sgdma_tx_csr_translator_avalon_anti_slave_0_read                                                      : std_logic;                      -- sgdma_tx_csr_translator:av_read -> sgdma_tx:csr_read
	signal sgdma_tx_csr_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(31 downto 0);  -- sgdma_tx:csr_readdata -> sgdma_tx_csr_translator:av_readdata
	signal sgdma_rx_csr_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(31 downto 0);  -- sgdma_rx_csr_translator:av_writedata -> sgdma_rx:csr_writedata
	signal sgdma_rx_csr_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(3 downto 0);   -- sgdma_rx_csr_translator:av_address -> sgdma_rx:csr_address
	signal sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect                                                : std_logic;                      -- sgdma_rx_csr_translator:av_chipselect -> sgdma_rx:csr_chipselect
	signal sgdma_rx_csr_translator_avalon_anti_slave_0_write                                                     : std_logic;                      -- sgdma_rx_csr_translator:av_write -> sgdma_rx:csr_write
	signal sgdma_rx_csr_translator_avalon_anti_slave_0_read                                                      : std_logic;                      -- sgdma_rx_csr_translator:av_read -> sgdma_rx:csr_read
	signal sgdma_rx_csr_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(31 downto 0);  -- sgdma_rx:csr_readdata -> sgdma_rx_csr_translator:av_readdata
	signal cpu_to_flash_ccb_m0_burstcount                                                                        : std_logic_vector(0 downto 0);   -- cpu_to_flash_ccb:m0_burstcount -> cpu_to_flash_ccb_m0_translator:av_burstcount
	signal cpu_to_flash_ccb_m0_waitrequest                                                                       : std_logic;                      -- cpu_to_flash_ccb_m0_translator:av_waitrequest -> cpu_to_flash_ccb:m0_waitrequest
	signal cpu_to_flash_ccb_m0_address                                                                           : std_logic_vector(27 downto 0);  -- cpu_to_flash_ccb:m0_address -> cpu_to_flash_ccb_m0_translator:av_address
	signal cpu_to_flash_ccb_m0_writedata                                                                         : std_logic_vector(31 downto 0);  -- cpu_to_flash_ccb:m0_writedata -> cpu_to_flash_ccb_m0_translator:av_writedata
	signal cpu_to_flash_ccb_m0_write                                                                             : std_logic;                      -- cpu_to_flash_ccb:m0_write -> cpu_to_flash_ccb_m0_translator:av_write
	signal cpu_to_flash_ccb_m0_read                                                                              : std_logic;                      -- cpu_to_flash_ccb:m0_read -> cpu_to_flash_ccb_m0_translator:av_read
	signal cpu_to_flash_ccb_m0_readdata                                                                          : std_logic_vector(31 downto 0);  -- cpu_to_flash_ccb_m0_translator:av_readdata -> cpu_to_flash_ccb:m0_readdata
	signal cpu_to_flash_ccb_m0_debugaccess                                                                       : std_logic;                      -- cpu_to_flash_ccb:m0_debugaccess -> cpu_to_flash_ccb_m0_translator:av_debugaccess
	signal cpu_to_flash_ccb_m0_byteenable                                                                        : std_logic_vector(3 downto 0);   -- cpu_to_flash_ccb:m0_byteenable -> cpu_to_flash_ccb_m0_translator:av_byteenable
	signal cpu_to_flash_ccb_m0_readdatavalid                                                                     : std_logic;                      -- cpu_to_flash_ccb_m0_translator:av_readdatavalid -> cpu_to_flash_ccb:m0_readdatavalid
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_waitrequest                           : std_logic;                      -- cfi_flash_ts_controller_fpga:uas_waitrequest -> cfi_flash_ts_controller_fpga_uas_translator:av_waitrequest
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_burstcount                            : std_logic_vector(1 downto 0);   -- cfi_flash_ts_controller_fpga_uas_translator:av_burstcount -> cfi_flash_ts_controller_fpga:uas_burstcount
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(15 downto 0);  -- cfi_flash_ts_controller_fpga_uas_translator:av_writedata -> cfi_flash_ts_controller_fpga:uas_writedata
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_address                               : std_logic_vector(26 downto 0);  -- cfi_flash_ts_controller_fpga_uas_translator:av_address -> cfi_flash_ts_controller_fpga:uas_address
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_lock                                  : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator:av_lock -> cfi_flash_ts_controller_fpga:uas_lock
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_write                                 : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator:av_write -> cfi_flash_ts_controller_fpga:uas_write
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_read                                  : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator:av_read -> cfi_flash_ts_controller_fpga:uas_read
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(15 downto 0);  -- cfi_flash_ts_controller_fpga:uas_readdata -> cfi_flash_ts_controller_fpga_uas_translator:av_readdata
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_debugaccess                           : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator:av_debugaccess -> cfi_flash_ts_controller_fpga:uas_debugaccess
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_readdatavalid                         : std_logic;                      -- cfi_flash_ts_controller_fpga:uas_readdatavalid -> cfi_flash_ts_controller_fpga_uas_translator:av_readdatavalid
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_byteenable                            : std_logic_vector(1 downto 0);   -- cfi_flash_ts_controller_fpga_uas_translator:av_byteenable -> cfi_flash_ts_controller_fpga:uas_byteenable
	signal cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_waitrequest                                : std_logic;                      -- cfi_flash_ts_controller:uas_waitrequest -> cfi_flash_ts_controller_uas_translator:av_waitrequest
	signal cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_burstcount                                 : std_logic_vector(1 downto 0);   -- cfi_flash_ts_controller_uas_translator:av_burstcount -> cfi_flash_ts_controller:uas_burstcount
	signal cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_writedata                                  : std_logic_vector(15 downto 0);  -- cfi_flash_ts_controller_uas_translator:av_writedata -> cfi_flash_ts_controller:uas_writedata
	signal cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_address                                    : std_logic_vector(26 downto 0);  -- cfi_flash_ts_controller_uas_translator:av_address -> cfi_flash_ts_controller:uas_address
	signal cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_lock                                       : std_logic;                      -- cfi_flash_ts_controller_uas_translator:av_lock -> cfi_flash_ts_controller:uas_lock
	signal cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_write                                      : std_logic;                      -- cfi_flash_ts_controller_uas_translator:av_write -> cfi_flash_ts_controller:uas_write
	signal cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_read                                       : std_logic;                      -- cfi_flash_ts_controller_uas_translator:av_read -> cfi_flash_ts_controller:uas_read
	signal cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_readdata                                   : std_logic_vector(15 downto 0);  -- cfi_flash_ts_controller:uas_readdata -> cfi_flash_ts_controller_uas_translator:av_readdata
	signal cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_debugaccess                                : std_logic;                      -- cfi_flash_ts_controller_uas_translator:av_debugaccess -> cfi_flash_ts_controller:uas_debugaccess
	signal cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_readdatavalid                              : std_logic;                      -- cfi_flash_ts_controller:uas_readdatavalid -> cfi_flash_ts_controller_uas_translator:av_readdatavalid
	signal cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_byteenable                                 : std_logic_vector(1 downto 0);   -- cfi_flash_ts_controller_uas_translator:av_byteenable -> cfi_flash_ts_controller:uas_byteenable
	signal sgdma_tx_m_read_waitrequest                                                                           : std_logic;                      -- sgdma_tx_m_read_translator:av_waitrequest -> sgdma_tx:m_read_waitrequest
	signal sgdma_tx_m_read_address                                                                               : std_logic_vector(31 downto 0);  -- sgdma_tx:m_read_address -> sgdma_tx_m_read_translator:av_address
	signal sgdma_tx_m_read_read                                                                                  : std_logic;                      -- sgdma_tx:m_read_read -> sgdma_tx_m_read_translator:av_read
	signal sgdma_tx_m_read_readdata                                                                              : std_logic_vector(31 downto 0);  -- sgdma_tx_m_read_translator:av_readdata -> sgdma_tx:m_read_readdata
	signal sgdma_tx_m_read_readdatavalid                                                                         : std_logic;                      -- sgdma_tx_m_read_translator:av_readdatavalid -> sgdma_tx:m_read_readdatavalid
	signal sgdma_rx_m_write_waitrequest                                                                          : std_logic;                      -- sgdma_rx_m_write_translator:av_waitrequest -> sgdma_rx:m_write_waitrequest
	signal sgdma_rx_m_write_writedata                                                                            : std_logic_vector(31 downto 0);  -- sgdma_rx:m_write_writedata -> sgdma_rx_m_write_translator:av_writedata
	signal sgdma_rx_m_write_address                                                                              : std_logic_vector(31 downto 0);  -- sgdma_rx:m_write_address -> sgdma_rx_m_write_translator:av_address
	signal sgdma_rx_m_write_write                                                                                : std_logic;                      -- sgdma_rx:m_write_write -> sgdma_rx_m_write_translator:av_write
	signal sgdma_rx_m_write_byteenable                                                                           : std_logic_vector(3 downto 0);   -- sgdma_rx:m_write_byteenable -> sgdma_rx_m_write_translator:av_byteenable
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_waitrequest                                    : std_logic;                      -- tse_dma_to_sdram_ccb:s0_waitrequest -> tse_dma_to_sdram_ccb_s0_translator:av_waitrequest
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_burstcount                                     : std_logic_vector(0 downto 0);   -- tse_dma_to_sdram_ccb_s0_translator:av_burstcount -> tse_dma_to_sdram_ccb:s0_burstcount
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_writedata                                      : std_logic_vector(31 downto 0);  -- tse_dma_to_sdram_ccb_s0_translator:av_writedata -> tse_dma_to_sdram_ccb:s0_writedata
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_address                                        : std_logic_vector(26 downto 0);  -- tse_dma_to_sdram_ccb_s0_translator:av_address -> tse_dma_to_sdram_ccb:s0_address
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_write                                          : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator:av_write -> tse_dma_to_sdram_ccb:s0_write
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_read                                           : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator:av_read -> tse_dma_to_sdram_ccb:s0_read
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_readdata                                       : std_logic_vector(31 downto 0);  -- tse_dma_to_sdram_ccb:s0_readdata -> tse_dma_to_sdram_ccb_s0_translator:av_readdata
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_debugaccess                                    : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator:av_debugaccess -> tse_dma_to_sdram_ccb:s0_debugaccess
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_readdatavalid                                  : std_logic;                      -- tse_dma_to_sdram_ccb:s0_readdatavalid -> tse_dma_to_sdram_ccb_s0_translator:av_readdatavalid
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_byteenable                                     : std_logic_vector(3 downto 0);   -- tse_dma_to_sdram_ccb_s0_translator:av_byteenable -> tse_dma_to_sdram_ccb:s0_byteenable
	signal tse_dma_to_sdram_ccb_m0_burstcount                                                                    : std_logic_vector(0 downto 0);   -- tse_dma_to_sdram_ccb:m0_burstcount -> tse_dma_to_sdram_ccb_m0_translator:av_burstcount
	signal tse_dma_to_sdram_ccb_m0_waitrequest                                                                   : std_logic;                      -- tse_dma_to_sdram_ccb_m0_translator:av_waitrequest -> tse_dma_to_sdram_ccb:m0_waitrequest
	signal tse_dma_to_sdram_ccb_m0_address                                                                       : std_logic_vector(26 downto 0);  -- tse_dma_to_sdram_ccb:m0_address -> tse_dma_to_sdram_ccb_m0_translator:av_address
	signal tse_dma_to_sdram_ccb_m0_writedata                                                                     : std_logic_vector(31 downto 0);  -- tse_dma_to_sdram_ccb:m0_writedata -> tse_dma_to_sdram_ccb_m0_translator:av_writedata
	signal tse_dma_to_sdram_ccb_m0_write                                                                         : std_logic;                      -- tse_dma_to_sdram_ccb:m0_write -> tse_dma_to_sdram_ccb_m0_translator:av_write
	signal tse_dma_to_sdram_ccb_m0_read                                                                          : std_logic;                      -- tse_dma_to_sdram_ccb:m0_read -> tse_dma_to_sdram_ccb_m0_translator:av_read
	signal tse_dma_to_sdram_ccb_m0_readdata                                                                      : std_logic_vector(31 downto 0);  -- tse_dma_to_sdram_ccb_m0_translator:av_readdata -> tse_dma_to_sdram_ccb:m0_readdata
	signal tse_dma_to_sdram_ccb_m0_debugaccess                                                                   : std_logic;                      -- tse_dma_to_sdram_ccb:m0_debugaccess -> tse_dma_to_sdram_ccb_m0_translator:av_debugaccess
	signal tse_dma_to_sdram_ccb_m0_byteenable                                                                    : std_logic_vector(3 downto 0);   -- tse_dma_to_sdram_ccb:m0_byteenable -> tse_dma_to_sdram_ccb_m0_translator:av_byteenable
	signal tse_dma_to_sdram_ccb_m0_readdatavalid                                                                 : std_logic;                      -- tse_dma_to_sdram_ccb_m0_translator:av_readdatavalid -> tse_dma_to_sdram_ccb:m0_readdatavalid
	signal cpu_to_sdram_pb_m0_burstcount                                                                         : std_logic_vector(0 downto 0);   -- cpu_to_sdram_pb:m0_burstcount -> cpu_to_sdram_pb_m0_translator:av_burstcount
	signal cpu_to_sdram_pb_m0_waitrequest                                                                        : std_logic;                      -- cpu_to_sdram_pb_m0_translator:av_waitrequest -> cpu_to_sdram_pb:m0_waitrequest
	signal cpu_to_sdram_pb_m0_address                                                                            : std_logic_vector(26 downto 0);  -- cpu_to_sdram_pb:m0_address -> cpu_to_sdram_pb_m0_translator:av_address
	signal cpu_to_sdram_pb_m0_writedata                                                                          : std_logic_vector(31 downto 0);  -- cpu_to_sdram_pb:m0_writedata -> cpu_to_sdram_pb_m0_translator:av_writedata
	signal cpu_to_sdram_pb_m0_write                                                                              : std_logic;                      -- cpu_to_sdram_pb:m0_write -> cpu_to_sdram_pb_m0_translator:av_write
	signal cpu_to_sdram_pb_m0_read                                                                               : std_logic;                      -- cpu_to_sdram_pb:m0_read -> cpu_to_sdram_pb_m0_translator:av_read
	signal cpu_to_sdram_pb_m0_readdata                                                                           : std_logic_vector(31 downto 0);  -- cpu_to_sdram_pb_m0_translator:av_readdata -> cpu_to_sdram_pb:m0_readdata
	signal cpu_to_sdram_pb_m0_debugaccess                                                                        : std_logic;                      -- cpu_to_sdram_pb:m0_debugaccess -> cpu_to_sdram_pb_m0_translator:av_debugaccess
	signal cpu_to_sdram_pb_m0_byteenable                                                                         : std_logic_vector(3 downto 0);   -- cpu_to_sdram_pb:m0_byteenable -> cpu_to_sdram_pb_m0_translator:av_byteenable
	signal cpu_to_sdram_pb_m0_readdatavalid                                                                      : std_logic;                      -- cpu_to_sdram_pb_m0_translator:av_readdatavalid -> cpu_to_sdram_pb:m0_readdatavalid
	signal sdram_0_avl_waitrequest                                                                               : std_logic;                      -- sdram_0:avl_ready -> sdram_0_avl_waitrequest:in
	signal sdram_0_avl_translator_avalon_anti_slave_0_burstcount                                                 : std_logic_vector(2 downto 0);   -- sdram_0_avl_translator:av_burstcount -> sdram_0:avl_size
	signal sdram_0_avl_translator_avalon_anti_slave_0_writedata                                                  : std_logic_vector(63 downto 0);  -- sdram_0_avl_translator:av_writedata -> sdram_0:avl_wdata
	signal sdram_0_avl_translator_avalon_anti_slave_0_address                                                    : std_logic_vector(23 downto 0);  -- sdram_0_avl_translator:av_address -> sdram_0:avl_addr
	signal sdram_0_avl_translator_avalon_anti_slave_0_write                                                      : std_logic;                      -- sdram_0_avl_translator:av_write -> sdram_0:avl_write_req
	signal sdram_0_avl_translator_avalon_anti_slave_0_beginbursttransfer                                         : std_logic;                      -- sdram_0_avl_translator:av_beginbursttransfer -> sdram_0:avl_burstbegin
	signal sdram_0_avl_translator_avalon_anti_slave_0_read                                                       : std_logic;                      -- sdram_0_avl_translator:av_read -> sdram_0:avl_read_req
	signal sdram_0_avl_translator_avalon_anti_slave_0_readdata                                                   : std_logic_vector(63 downto 0);  -- sdram_0:avl_rdata -> sdram_0_avl_translator:av_readdata
	signal sdram_0_avl_translator_avalon_anti_slave_0_readdatavalid                                              : std_logic;                      -- sdram_0:avl_rdata_valid -> sdram_0_avl_translator:av_readdatavalid
	signal sdram_0_avl_translator_avalon_anti_slave_0_byteenable                                                 : std_logic_vector(7 downto 0);   -- sdram_0_avl_translator:av_byteenable -> sdram_0:avl_be
	signal linux_cpu_tightly_coupled_data_master_0_waitrequest                                                   : std_logic;                      -- linux_cpu_tightly_coupled_data_master_0_translator:av_waitrequest -> linux_cpu:dcm0_waitrequest
	signal linux_cpu_tightly_coupled_data_master_0_writedata                                                     : std_logic_vector(31 downto 0);  -- linux_cpu:dcm0_writedata -> linux_cpu_tightly_coupled_data_master_0_translator:av_writedata
	signal linux_cpu_tightly_coupled_data_master_0_address                                                       : std_logic_vector(28 downto 0);  -- linux_cpu:dcm0_address -> linux_cpu_tightly_coupled_data_master_0_translator:av_address
	signal linux_cpu_tightly_coupled_data_master_0_clken                                                         : std_logic;                      -- linux_cpu:dcm0_clken -> linux_cpu_tightly_coupled_data_master_0_translator:av_clken
	signal linux_cpu_tightly_coupled_data_master_0_write                                                         : std_logic;                      -- linux_cpu:dcm0_write -> linux_cpu_tightly_coupled_data_master_0_translator:av_write
	signal linux_cpu_tightly_coupled_data_master_0_read                                                          : std_logic;                      -- linux_cpu:dcm0_read -> linux_cpu_tightly_coupled_data_master_0_translator:av_read
	signal linux_cpu_tightly_coupled_data_master_0_readdata                                                      : std_logic_vector(31 downto 0);  -- linux_cpu_tightly_coupled_data_master_0_translator:av_readdata -> linux_cpu:dcm0_readdata
	signal linux_cpu_tightly_coupled_data_master_0_byteenable                                                    : std_logic_vector(3 downto 0);   -- linux_cpu:dcm0_byteenable -> linux_cpu_tightly_coupled_data_master_0_translator:av_byteenable
	signal linux_cpu_tightly_coupled_data_master_0_readdatavalid                                                 : std_logic;                      -- linux_cpu_tightly_coupled_data_master_0_translator:av_readdatavalid -> linux_cpu:dcm0_readdatavalid
	signal linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_waitrequest              : std_logic;                      -- tlb_miss_ram_1k_s1_translator:uav_waitrequest -> linux_cpu_tightly_coupled_data_master_0_translator:uav_waitrequest
	signal linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_burstcount               : std_logic_vector(2 downto 0);   -- linux_cpu_tightly_coupled_data_master_0_translator:uav_burstcount -> tlb_miss_ram_1k_s1_translator:uav_burstcount
	signal linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_writedata                : std_logic_vector(31 downto 0);  -- linux_cpu_tightly_coupled_data_master_0_translator:uav_writedata -> tlb_miss_ram_1k_s1_translator:uav_writedata
	signal linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_address                  : std_logic_vector(28 downto 0);  -- linux_cpu_tightly_coupled_data_master_0_translator:uav_address -> tlb_miss_ram_1k_s1_translator:uav_address
	signal linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_clken                    : std_logic;                      -- linux_cpu_tightly_coupled_data_master_0_translator:uav_clken -> tlb_miss_ram_1k_s1_translator:uav_clken
	signal linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_lock                     : std_logic;                      -- linux_cpu_tightly_coupled_data_master_0_translator:uav_lock -> tlb_miss_ram_1k_s1_translator:uav_lock
	signal linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_write                    : std_logic;                      -- linux_cpu_tightly_coupled_data_master_0_translator:uav_write -> tlb_miss_ram_1k_s1_translator:uav_write
	signal linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_read                     : std_logic;                      -- linux_cpu_tightly_coupled_data_master_0_translator:uav_read -> tlb_miss_ram_1k_s1_translator:uav_read
	signal linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_readdata                 : std_logic_vector(31 downto 0);  -- tlb_miss_ram_1k_s1_translator:uav_readdata -> linux_cpu_tightly_coupled_data_master_0_translator:uav_readdata
	signal linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_debugaccess              : std_logic;                      -- linux_cpu_tightly_coupled_data_master_0_translator:uav_debugaccess -> tlb_miss_ram_1k_s1_translator:uav_debugaccess
	signal linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_byteenable               : std_logic_vector(3 downto 0);   -- linux_cpu_tightly_coupled_data_master_0_translator:uav_byteenable -> tlb_miss_ram_1k_s1_translator:uav_byteenable
	signal linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_readdatavalid            : std_logic;                      -- tlb_miss_ram_1k_s1_translator:uav_readdatavalid -> linux_cpu_tightly_coupled_data_master_0_translator:uav_readdatavalid
	signal tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_writedata                                           : std_logic_vector(31 downto 0);  -- tlb_miss_ram_1k_s1_translator:av_writedata -> tlb_miss_ram_1k:writedata
	signal tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_address                                             : std_logic_vector(7 downto 0);   -- tlb_miss_ram_1k_s1_translator:av_address -> tlb_miss_ram_1k:address
	signal tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_chipselect                                          : std_logic;                      -- tlb_miss_ram_1k_s1_translator:av_chipselect -> tlb_miss_ram_1k:chipselect
	signal tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_clken                                               : std_logic;                      -- tlb_miss_ram_1k_s1_translator:av_clken -> tlb_miss_ram_1k:clken
	signal tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_write                                               : std_logic;                      -- tlb_miss_ram_1k_s1_translator:av_write -> tlb_miss_ram_1k:write
	signal tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_readdata                                            : std_logic_vector(31 downto 0);  -- tlb_miss_ram_1k:readdata -> tlb_miss_ram_1k_s1_translator:av_readdata
	signal tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_byteenable                                          : std_logic_vector(3 downto 0);   -- tlb_miss_ram_1k_s1_translator:av_byteenable -> tlb_miss_ram_1k:byteenable
	signal linux_cpu_tightly_coupled_instruction_master_0_waitrequest                                            : std_logic;                      -- linux_cpu_tightly_coupled_instruction_master_0_translator:av_waitrequest -> linux_cpu:icm0_waitrequest
	signal linux_cpu_tightly_coupled_instruction_master_0_address                                                : std_logic_vector(28 downto 0);  -- linux_cpu:icm0_address -> linux_cpu_tightly_coupled_instruction_master_0_translator:av_address
	signal linux_cpu_tightly_coupled_instruction_master_0_clken                                                  : std_logic;                      -- linux_cpu:icm0_clken -> linux_cpu_tightly_coupled_instruction_master_0_translator:av_clken
	signal linux_cpu_tightly_coupled_instruction_master_0_read                                                   : std_logic;                      -- linux_cpu:icm0_read -> linux_cpu_tightly_coupled_instruction_master_0_translator:av_read
	signal linux_cpu_tightly_coupled_instruction_master_0_readdata                                               : std_logic_vector(31 downto 0);  -- linux_cpu_tightly_coupled_instruction_master_0_translator:av_readdata -> linux_cpu:icm0_readdata
	signal linux_cpu_tightly_coupled_instruction_master_0_readdatavalid                                          : std_logic;                      -- linux_cpu_tightly_coupled_instruction_master_0_translator:av_readdatavalid -> linux_cpu:icm0_readdatavalid
	signal linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_waitrequest       : std_logic;                      -- tlb_miss_ram_1k_s2_translator:uav_waitrequest -> linux_cpu_tightly_coupled_instruction_master_0_translator:uav_waitrequest
	signal linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_burstcount        : std_logic_vector(2 downto 0);   -- linux_cpu_tightly_coupled_instruction_master_0_translator:uav_burstcount -> tlb_miss_ram_1k_s2_translator:uav_burstcount
	signal linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_writedata         : std_logic_vector(31 downto 0);  -- linux_cpu_tightly_coupled_instruction_master_0_translator:uav_writedata -> tlb_miss_ram_1k_s2_translator:uav_writedata
	signal linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_address           : std_logic_vector(28 downto 0);  -- linux_cpu_tightly_coupled_instruction_master_0_translator:uav_address -> tlb_miss_ram_1k_s2_translator:uav_address
	signal linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_clken             : std_logic;                      -- linux_cpu_tightly_coupled_instruction_master_0_translator:uav_clken -> tlb_miss_ram_1k_s2_translator:uav_clken
	signal linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_lock              : std_logic;                      -- linux_cpu_tightly_coupled_instruction_master_0_translator:uav_lock -> tlb_miss_ram_1k_s2_translator:uav_lock
	signal linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_write             : std_logic;                      -- linux_cpu_tightly_coupled_instruction_master_0_translator:uav_write -> tlb_miss_ram_1k_s2_translator:uav_write
	signal linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_read              : std_logic;                      -- linux_cpu_tightly_coupled_instruction_master_0_translator:uav_read -> tlb_miss_ram_1k_s2_translator:uav_read
	signal linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_readdata          : std_logic_vector(31 downto 0);  -- tlb_miss_ram_1k_s2_translator:uav_readdata -> linux_cpu_tightly_coupled_instruction_master_0_translator:uav_readdata
	signal linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_debugaccess       : std_logic;                      -- linux_cpu_tightly_coupled_instruction_master_0_translator:uav_debugaccess -> tlb_miss_ram_1k_s2_translator:uav_debugaccess
	signal linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_byteenable        : std_logic_vector(3 downto 0);   -- linux_cpu_tightly_coupled_instruction_master_0_translator:uav_byteenable -> tlb_miss_ram_1k_s2_translator:uav_byteenable
	signal linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_readdatavalid     : std_logic;                      -- tlb_miss_ram_1k_s2_translator:uav_readdatavalid -> linux_cpu_tightly_coupled_instruction_master_0_translator:uav_readdatavalid
	signal tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_writedata                                           : std_logic_vector(31 downto 0);  -- tlb_miss_ram_1k_s2_translator:av_writedata -> tlb_miss_ram_1k:writedata2
	signal tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_address                                             : std_logic_vector(7 downto 0);   -- tlb_miss_ram_1k_s2_translator:av_address -> tlb_miss_ram_1k:address2
	signal tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_chipselect                                          : std_logic;                      -- tlb_miss_ram_1k_s2_translator:av_chipselect -> tlb_miss_ram_1k:chipselect2
	signal tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_clken                                               : std_logic;                      -- tlb_miss_ram_1k_s2_translator:av_clken -> tlb_miss_ram_1k:clken2
	signal tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_write                                               : std_logic;                      -- tlb_miss_ram_1k_s2_translator:av_write -> tlb_miss_ram_1k:write2
	signal tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_readdata                                            : std_logic_vector(31 downto 0);  -- tlb_miss_ram_1k:readdata2 -> tlb_miss_ram_1k_s2_translator:av_readdata
	signal tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_byteenable                                          : std_logic_vector(3 downto 0);   -- tlb_miss_ram_1k_s2_translator:av_byteenable -> tlb_miss_ram_1k:byteenable2
	signal linux_cpu_data_master_translator_avalon_universal_master_0_waitrequest                                : std_logic;                      -- linux_cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> linux_cpu_data_master_translator:uav_waitrequest
	signal linux_cpu_data_master_translator_avalon_universal_master_0_burstcount                                 : std_logic_vector(2 downto 0);   -- linux_cpu_data_master_translator:uav_burstcount -> linux_cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal linux_cpu_data_master_translator_avalon_universal_master_0_writedata                                  : std_logic_vector(31 downto 0);  -- linux_cpu_data_master_translator:uav_writedata -> linux_cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal linux_cpu_data_master_translator_avalon_universal_master_0_address                                    : std_logic_vector(28 downto 0);  -- linux_cpu_data_master_translator:uav_address -> linux_cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	signal linux_cpu_data_master_translator_avalon_universal_master_0_lock                                       : std_logic;                      -- linux_cpu_data_master_translator:uav_lock -> linux_cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal linux_cpu_data_master_translator_avalon_universal_master_0_write                                      : std_logic;                      -- linux_cpu_data_master_translator:uav_write -> linux_cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	signal linux_cpu_data_master_translator_avalon_universal_master_0_read                                       : std_logic;                      -- linux_cpu_data_master_translator:uav_read -> linux_cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	signal linux_cpu_data_master_translator_avalon_universal_master_0_readdata                                   : std_logic_vector(31 downto 0);  -- linux_cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> linux_cpu_data_master_translator:uav_readdata
	signal linux_cpu_data_master_translator_avalon_universal_master_0_debugaccess                                : std_logic;                      -- linux_cpu_data_master_translator:uav_debugaccess -> linux_cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal linux_cpu_data_master_translator_avalon_universal_master_0_byteenable                                 : std_logic_vector(3 downto 0);   -- linux_cpu_data_master_translator:uav_byteenable -> linux_cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal linux_cpu_data_master_translator_avalon_universal_master_0_readdatavalid                              : std_logic;                      -- linux_cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> linux_cpu_data_master_translator:uav_readdatavalid
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_waitrequest                         : std_logic;                      -- linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> linux_cpu_instruction_master_translator:uav_waitrequest
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_burstcount                          : std_logic_vector(2 downto 0);   -- linux_cpu_instruction_master_translator:uav_burstcount -> linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_writedata                           : std_logic_vector(31 downto 0);  -- linux_cpu_instruction_master_translator:uav_writedata -> linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_address                             : std_logic_vector(28 downto 0);  -- linux_cpu_instruction_master_translator:uav_address -> linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_lock                                : std_logic;                      -- linux_cpu_instruction_master_translator:uav_lock -> linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_write                               : std_logic;                      -- linux_cpu_instruction_master_translator:uav_write -> linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_read                                : std_logic;                      -- linux_cpu_instruction_master_translator:uav_read -> linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_readdata                            : std_logic_vector(31 downto 0);  -- linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> linux_cpu_instruction_master_translator:uav_readdata
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_debugaccess                         : std_logic;                      -- linux_cpu_instruction_master_translator:uav_debugaccess -> linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_byteenable                          : std_logic_vector(3 downto 0);   -- linux_cpu_instruction_master_translator:uav_byteenable -> linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid                       : std_logic;                      -- linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> linux_cpu_instruction_master_translator:uav_readdatavalid
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest                  : std_logic;                      -- linux_cpu_jtag_debug_module_translator:uav_waitrequest -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount                   : std_logic_vector(2 downto 0);   -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> linux_cpu_jtag_debug_module_translator:uav_burstcount
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata                    : std_logic_vector(31 downto 0);  -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> linux_cpu_jtag_debug_module_translator:uav_writedata
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                      : std_logic_vector(28 downto 0);  -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> linux_cpu_jtag_debug_module_translator:uav_address
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                        : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> linux_cpu_jtag_debug_module_translator:uav_write
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                         : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> linux_cpu_jtag_debug_module_translator:uav_lock
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                         : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> linux_cpu_jtag_debug_module_translator:uav_read
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                     : std_logic_vector(31 downto 0);  -- linux_cpu_jtag_debug_module_translator:uav_readdata -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid                : std_logic;                      -- linux_cpu_jtag_debug_module_translator:uav_readdatavalid -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess                  : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> linux_cpu_jtag_debug_module_translator:uav_debugaccess
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable                   : std_logic_vector(3 downto 0);   -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> linux_cpu_jtag_debug_module_translator:uav_byteenable
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket           : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid                 : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket         : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data                  : std_logic_vector(100 downto 0); -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready                 : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket        : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid              : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket      : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data               : std_logic_vector(100 downto 0); -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready              : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid            : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data             : std_logic_vector(33 downto 0);  -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready            : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest                          : std_logic;                      -- cpu_to_flash_ccb_s0_translator:uav_waitrequest -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount                           : std_logic_vector(2 downto 0);   -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_to_flash_ccb_s0_translator:uav_burstcount
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_writedata                            : std_logic_vector(31 downto 0);  -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_to_flash_ccb_s0_translator:uav_writedata
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_address                              : std_logic_vector(28 downto 0);  -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:m0_address -> cpu_to_flash_ccb_s0_translator:uav_address
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_write                                : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:m0_write -> cpu_to_flash_ccb_s0_translator:uav_write
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_lock                                 : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_to_flash_ccb_s0_translator:uav_lock
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_read                                 : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:m0_read -> cpu_to_flash_ccb_s0_translator:uav_read
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdata                             : std_logic_vector(31 downto 0);  -- cpu_to_flash_ccb_s0_translator:uav_readdata -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                        : std_logic;                      -- cpu_to_flash_ccb_s0_translator:uav_readdatavalid -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess                          : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_to_flash_ccb_s0_translator:uav_debugaccess
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable                           : std_logic_vector(3 downto 0);   -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_to_flash_ccb_s0_translator:uav_byteenable
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                   : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid                         : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                 : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_data                          : std_logic_vector(100 downto 0); -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready                         : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                      : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket              : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                       : std_logic_vector(100 downto 0); -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                      : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                    : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                     : std_logic_vector(33 downto 0);  -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                    : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest                    : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator:uav_waitrequest -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount                     : std_logic_vector(2 downto 0);   -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_to_peripherals_ccb_s0_translator:uav_burstcount
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_writedata                      : std_logic_vector(31 downto 0);  -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_to_peripherals_ccb_s0_translator:uav_writedata
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_address                        : std_logic_vector(28 downto 0);  -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:m0_address -> cpu_to_peripherals_ccb_s0_translator:uav_address
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_write                          : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:m0_write -> cpu_to_peripherals_ccb_s0_translator:uav_write
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_lock                           : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_to_peripherals_ccb_s0_translator:uav_lock
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_read                           : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:m0_read -> cpu_to_peripherals_ccb_s0_translator:uav_read
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdata                       : std_logic_vector(31 downto 0);  -- cpu_to_peripherals_ccb_s0_translator:uav_readdata -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                  : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator:uav_readdatavalid -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess                    : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_to_peripherals_ccb_s0_translator:uav_debugaccess
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable                     : std_logic_vector(3 downto 0);   -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_to_peripherals_ccb_s0_translator:uav_byteenable
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket             : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid                   : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket           : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_data                    : std_logic_vector(100 downto 0); -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready                   : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket          : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket        : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                 : std_logic_vector(100 downto 0); -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid              : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data               : std_logic_vector(33 downto 0);  -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready              : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest                           : std_logic;                      -- cpu_to_sdram_pb_s0_translator:uav_waitrequest -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount                            : std_logic_vector(2 downto 0);   -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_to_sdram_pb_s0_translator:uav_burstcount
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_writedata                             : std_logic_vector(31 downto 0);  -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_to_sdram_pb_s0_translator:uav_writedata
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_address                               : std_logic_vector(28 downto 0);  -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:m0_address -> cpu_to_sdram_pb_s0_translator:uav_address
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_write                                 : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:m0_write -> cpu_to_sdram_pb_s0_translator:uav_write
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_lock                                  : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_to_sdram_pb_s0_translator:uav_lock
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_read                                  : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:m0_read -> cpu_to_sdram_pb_s0_translator:uav_read
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_readdata                              : std_logic_vector(31 downto 0);  -- cpu_to_sdram_pb_s0_translator:uav_readdata -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                         : std_logic;                      -- cpu_to_sdram_pb_s0_translator:uav_readdatavalid -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess                           : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_to_sdram_pb_s0_translator:uav_debugaccess
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable                            : std_logic_vector(3 downto 0);   -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_to_sdram_pb_s0_translator:uav_byteenable
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                    : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid                          : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                  : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rf_source_data                           : std_logic_vector(100 downto 0); -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready                          : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                 : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                       : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket               : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                        : std_logic_vector(100 downto 0); -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                       : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                     : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                      : std_logic_vector(33 downto 0);  -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                     : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest                            : std_logic;                      -- sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_descriptor_write_translator:uav_waitrequest
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount                             : std_logic_vector(2 downto 0);   -- sgdma_tx_descriptor_write_translator:uav_burstcount -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_burstcount
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata                              : std_logic_vector(31 downto 0);  -- sgdma_tx_descriptor_write_translator:uav_writedata -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_writedata
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address                                : std_logic_vector(31 downto 0);  -- sgdma_tx_descriptor_write_translator:uav_address -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_address
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock                                   : std_logic;                      -- sgdma_tx_descriptor_write_translator:uav_lock -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_lock
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write                                  : std_logic;                      -- sgdma_tx_descriptor_write_translator:uav_write -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_write
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read                                   : std_logic;                      -- sgdma_tx_descriptor_write_translator:uav_read -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_read
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata                               : std_logic_vector(31 downto 0);  -- sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_descriptor_write_translator:uav_readdata
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess                            : std_logic;                      -- sgdma_tx_descriptor_write_translator:uav_debugaccess -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_debugaccess
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable                             : std_logic_vector(3 downto 0);   -- sgdma_tx_descriptor_write_translator:uav_byteenable -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_byteenable
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid                          : std_logic;                      -- sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_descriptor_write_translator:uav_readdatavalid
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest                            : std_logic;                      -- sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_descriptor_write_translator:uav_waitrequest
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount                             : std_logic_vector(2 downto 0);   -- sgdma_rx_descriptor_write_translator:uav_burstcount -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_burstcount
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata                              : std_logic_vector(31 downto 0);  -- sgdma_rx_descriptor_write_translator:uav_writedata -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_writedata
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address                                : std_logic_vector(31 downto 0);  -- sgdma_rx_descriptor_write_translator:uav_address -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_address
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock                                   : std_logic;                      -- sgdma_rx_descriptor_write_translator:uav_lock -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_lock
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write                                  : std_logic;                      -- sgdma_rx_descriptor_write_translator:uav_write -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_write
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read                                   : std_logic;                      -- sgdma_rx_descriptor_write_translator:uav_read -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_read
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata                               : std_logic_vector(31 downto 0);  -- sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_descriptor_write_translator:uav_readdata
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess                            : std_logic;                      -- sgdma_rx_descriptor_write_translator:uav_debugaccess -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_debugaccess
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable                             : std_logic_vector(3 downto 0);   -- sgdma_rx_descriptor_write_translator:uav_byteenable -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_byteenable
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid                          : std_logic;                      -- sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_descriptor_write_translator:uav_readdatavalid
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest                             : std_logic;                      -- sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_descriptor_read_translator:uav_waitrequest
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount                              : std_logic_vector(2 downto 0);   -- sgdma_rx_descriptor_read_translator:uav_burstcount -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_burstcount
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata                               : std_logic_vector(31 downto 0);  -- sgdma_rx_descriptor_read_translator:uav_writedata -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_writedata
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address                                 : std_logic_vector(31 downto 0);  -- sgdma_rx_descriptor_read_translator:uav_address -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_address
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock                                    : std_logic;                      -- sgdma_rx_descriptor_read_translator:uav_lock -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_lock
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write                                   : std_logic;                      -- sgdma_rx_descriptor_read_translator:uav_write -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_write
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read                                    : std_logic;                      -- sgdma_rx_descriptor_read_translator:uav_read -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_read
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata                                : std_logic_vector(31 downto 0);  -- sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_descriptor_read_translator:uav_readdata
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess                             : std_logic;                      -- sgdma_rx_descriptor_read_translator:uav_debugaccess -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_debugaccess
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable                              : std_logic_vector(3 downto 0);   -- sgdma_rx_descriptor_read_translator:uav_byteenable -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_byteenable
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid                           : std_logic;                      -- sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_descriptor_read_translator:uav_readdatavalid
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest                             : std_logic;                      -- sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_descriptor_read_translator:uav_waitrequest
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount                              : std_logic_vector(2 downto 0);   -- sgdma_tx_descriptor_read_translator:uav_burstcount -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_burstcount
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata                               : std_logic_vector(31 downto 0);  -- sgdma_tx_descriptor_read_translator:uav_writedata -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_writedata
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address                                 : std_logic_vector(31 downto 0);  -- sgdma_tx_descriptor_read_translator:uav_address -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_address
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock                                    : std_logic;                      -- sgdma_tx_descriptor_read_translator:uav_lock -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_lock
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write                                   : std_logic;                      -- sgdma_tx_descriptor_read_translator:uav_write -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_write
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read                                    : std_logic;                      -- sgdma_tx_descriptor_read_translator:uav_read -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_read
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata                                : std_logic_vector(31 downto 0);  -- sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_descriptor_read_translator:uav_readdata
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess                             : std_logic;                      -- sgdma_tx_descriptor_read_translator:uav_debugaccess -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_debugaccess
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable                              : std_logic_vector(3 downto 0);   -- sgdma_tx_descriptor_read_translator:uav_byteenable -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_byteenable
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid                           : std_logic;                      -- sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_descriptor_read_translator:uav_readdatavalid
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest                     : std_logic;                      -- dma_to_descriptor_mem_s0_translator:uav_waitrequest -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_burstcount                      : std_logic_vector(2 downto 0);   -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> dma_to_descriptor_mem_s0_translator:uav_burstcount
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_writedata                       : std_logic_vector(31 downto 0);  -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> dma_to_descriptor_mem_s0_translator:uav_writedata
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_address                         : std_logic_vector(31 downto 0);  -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:m0_address -> dma_to_descriptor_mem_s0_translator:uav_address
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_write                           : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:m0_write -> dma_to_descriptor_mem_s0_translator:uav_write
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_lock                            : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:m0_lock -> dma_to_descriptor_mem_s0_translator:uav_lock
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_read                            : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:m0_read -> dma_to_descriptor_mem_s0_translator:uav_read
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_readdata                        : std_logic_vector(31 downto 0);  -- dma_to_descriptor_mem_s0_translator:uav_readdata -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                   : std_logic;                      -- dma_to_descriptor_mem_s0_translator:uav_readdatavalid -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess                     : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dma_to_descriptor_mem_s0_translator:uav_debugaccess
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_byteenable                      : std_logic_vector(3 downto 0);   -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> dma_to_descriptor_mem_s0_translator:uav_byteenable
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket              : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rf_source_valid                    : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket            : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rf_source_data                     : std_logic_vector(101 downto 0); -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rf_source_ready                    : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket           : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                 : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket         : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                  : std_logic_vector(101 downto 0); -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                 : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid               : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                : std_logic_vector(33 downto 0);  -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready               : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_waitrequest                             : std_logic;                      -- dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_to_descriptor_mem_m0_translator:uav_waitrequest
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_burstcount                              : std_logic_vector(2 downto 0);   -- dma_to_descriptor_mem_m0_translator:uav_burstcount -> dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:av_burstcount
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_writedata                               : std_logic_vector(31 downto 0);  -- dma_to_descriptor_mem_m0_translator:uav_writedata -> dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:av_writedata
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_address                                 : std_logic_vector(22 downto 0);  -- dma_to_descriptor_mem_m0_translator:uav_address -> dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:av_address
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_lock                                    : std_logic;                      -- dma_to_descriptor_mem_m0_translator:uav_lock -> dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:av_lock
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_write                                   : std_logic;                      -- dma_to_descriptor_mem_m0_translator:uav_write -> dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:av_write
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_read                                    : std_logic;                      -- dma_to_descriptor_mem_m0_translator:uav_read -> dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:av_read
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_readdata                                : std_logic_vector(31 downto 0);  -- dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:av_readdata -> dma_to_descriptor_mem_m0_translator:uav_readdata
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_debugaccess                             : std_logic;                      -- dma_to_descriptor_mem_m0_translator:uav_debugaccess -> dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_byteenable                              : std_logic_vector(3 downto 0);   -- dma_to_descriptor_mem_m0_translator:uav_byteenable -> dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:av_byteenable
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_readdatavalid                           : std_logic;                      -- dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_to_descriptor_mem_m0_translator:uav_readdatavalid
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_waitrequest                            : std_logic;                      -- cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_to_peripherals_ccb_m0_translator:uav_waitrequest
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_burstcount                             : std_logic_vector(2 downto 0);   -- cpu_to_peripherals_ccb_m0_translator:uav_burstcount -> cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_writedata                              : std_logic_vector(31 downto 0);  -- cpu_to_peripherals_ccb_m0_translator:uav_writedata -> cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_address                                : std_logic_vector(22 downto 0);  -- cpu_to_peripherals_ccb_m0_translator:uav_address -> cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:av_address
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_lock                                   : std_logic;                      -- cpu_to_peripherals_ccb_m0_translator:uav_lock -> cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_write                                  : std_logic;                      -- cpu_to_peripherals_ccb_m0_translator:uav_write -> cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:av_write
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_read                                   : std_logic;                      -- cpu_to_peripherals_ccb_m0_translator:uav_read -> cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:av_read
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_readdata                               : std_logic_vector(31 downto 0);  -- cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:av_readdata -> cpu_to_peripherals_ccb_m0_translator:uav_readdata
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_debugaccess                            : std_logic;                      -- cpu_to_peripherals_ccb_m0_translator:uav_debugaccess -> cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_byteenable                             : std_logic_vector(3 downto 0);   -- cpu_to_peripherals_ccb_m0_translator:uav_byteenable -> cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_readdatavalid                          : std_logic;                      -- cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_to_peripherals_ccb_m0_translator:uav_readdatavalid
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                         : std_logic;                      -- descriptor_memory_s1_translator:uav_waitrequest -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                          : std_logic_vector(2 downto 0);   -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> descriptor_memory_s1_translator:uav_burstcount
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata                           : std_logic_vector(31 downto 0);  -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> descriptor_memory_s1_translator:uav_writedata
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address                             : std_logic_vector(22 downto 0);  -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> descriptor_memory_s1_translator:uav_address
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write                               : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> descriptor_memory_s1_translator:uav_write
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock                                : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> descriptor_memory_s1_translator:uav_lock
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read                                : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> descriptor_memory_s1_translator:uav_read
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata                            : std_logic_vector(31 downto 0);  -- descriptor_memory_s1_translator:uav_readdata -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                       : std_logic;                      -- descriptor_memory_s1_translator:uav_readdatavalid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                         : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> descriptor_memory_s1_translator:uav_debugaccess
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                          : std_logic_vector(3 downto 0);   -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> descriptor_memory_s1_translator:uav_byteenable
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                  : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                        : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data                         : std_logic_vector(94 downto 0);  -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                        : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket               : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                     : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket             : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                      : std_logic_vector(94 downto 0);  -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                     : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                   : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                    : std_logic_vector(33 downto 0);  -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                   : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                  : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                   : std_logic_vector(2 downto 0);   -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                    : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                      : std_logic_vector(22 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                        : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                         : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                         : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                     : std_logic_vector(31 downto 0);  -- jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                  : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                   : std_logic_vector(3 downto 0);   -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket           : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                 : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket         : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data                  : std_logic_vector(94 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                 : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket        : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid              : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket      : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data               : std_logic_vector(94 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready              : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid            : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data             : std_logic_vector(33 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready            : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest                         : std_logic;                      -- tse_mac_control_port_translator:uav_waitrequest -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount                          : std_logic_vector(2 downto 0);   -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> tse_mac_control_port_translator:uav_burstcount
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata                           : std_logic_vector(31 downto 0);  -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> tse_mac_control_port_translator:uav_writedata
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address                             : std_logic_vector(22 downto 0);  -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_address -> tse_mac_control_port_translator:uav_address
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write                               : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_write -> tse_mac_control_port_translator:uav_write
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock                                : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> tse_mac_control_port_translator:uav_lock
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read                                : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_read -> tse_mac_control_port_translator:uav_read
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata                            : std_logic_vector(31 downto 0);  -- tse_mac_control_port_translator:uav_readdata -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid                       : std_logic;                      -- tse_mac_control_port_translator:uav_readdatavalid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess                         : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> tse_mac_control_port_translator:uav_debugaccess
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable                          : std_logic_vector(3 downto 0);   -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> tse_mac_control_port_translator:uav_byteenable
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                  : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid                        : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data                         : std_logic_vector(94 downto 0);  -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready                        : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket               : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                     : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket             : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                      : std_logic_vector(94 downto 0);  -- tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                     : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                   : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                    : std_logic_vector(33 downto 0);  -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                   : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                          : std_logic;                      -- sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                           : std_logic_vector(2 downto 0);   -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                            : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address                              : std_logic_vector(22 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write                                : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                                 : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read                                 : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                             : std_logic_vector(31 downto 0);  -- sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                        : std_logic;                      -- sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                          : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                           : std_logic_vector(3 downto 0);   -- sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                   : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                         : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                 : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                          : std_logic_vector(94 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                         : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                      : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket              : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                       : std_logic_vector(94 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                      : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                    : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                     : std_logic_vector(33 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                    : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                           : std_logic;                      -- linux_timer_1ms_s1_translator:uav_waitrequest -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                            : std_logic_vector(2 downto 0);   -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> linux_timer_1ms_s1_translator:uav_burstcount
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_writedata                             : std_logic_vector(31 downto 0);  -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> linux_timer_1ms_s1_translator:uav_writedata
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_address                               : std_logic_vector(22 downto 0);  -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:m0_address -> linux_timer_1ms_s1_translator:uav_address
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_write                                 : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:m0_write -> linux_timer_1ms_s1_translator:uav_write
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_lock                                  : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:m0_lock -> linux_timer_1ms_s1_translator:uav_lock
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_read                                  : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:m0_read -> linux_timer_1ms_s1_translator:uav_read
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_readdata                              : std_logic_vector(31 downto 0);  -- linux_timer_1ms_s1_translator:uav_readdata -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                         : std_logic;                      -- linux_timer_1ms_s1_translator:uav_readdatavalid -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                           : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> linux_timer_1ms_s1_translator:uav_debugaccess
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                            : std_logic_vector(3 downto 0);   -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> linux_timer_1ms_s1_translator:uav_byteenable
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                    : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                          : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                  : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rf_source_data                           : std_logic_vector(94 downto 0);  -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                          : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                 : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                       : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket               : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                        : std_logic_vector(94 downto 0);  -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                       : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                     : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                      : std_logic_vector(33 downto 0);  -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                     : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest                               : std_logic;                      -- gtp_regif_0_s0_translator:uav_waitrequest -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount                                : std_logic_vector(2 downto 0);   -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> gtp_regif_0_s0_translator:uav_burstcount
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata                                 : std_logic_vector(31 downto 0);  -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> gtp_regif_0_s0_translator:uav_writedata
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_address                                   : std_logic_vector(22 downto 0);  -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:m0_address -> gtp_regif_0_s0_translator:uav_address
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_write                                     : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:m0_write -> gtp_regif_0_s0_translator:uav_write
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_lock                                      : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:m0_lock -> gtp_regif_0_s0_translator:uav_lock
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_read                                      : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:m0_read -> gtp_regif_0_s0_translator:uav_read
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata                                  : std_logic_vector(31 downto 0);  -- gtp_regif_0_s0_translator:uav_readdata -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                             : std_logic;                      -- gtp_regif_0_s0_translator:uav_readdatavalid -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess                               : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> gtp_regif_0_s0_translator:uav_debugaccess
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable                                : std_logic_vector(3 downto 0);   -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> gtp_regif_0_s0_translator:uav_byteenable
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                        : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid                              : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                      : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data                               : std_logic_vector(94 downto 0);  -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready                              : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                     : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                           : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                   : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                            : std_logic_vector(94 downto 0);  -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                           : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                         : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                          : std_logic_vector(33 downto 0);  -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                         : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                      -- sgdma_tx_csr_translator:uav_waitrequest -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);   -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> sgdma_tx_csr_translator:uav_burstcount
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0);  -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> sgdma_tx_csr_translator:uav_writedata
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(22 downto 0);  -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_address -> sgdma_tx_csr_translator:uav_address
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_write -> sgdma_tx_csr_translator:uav_write
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_lock -> sgdma_tx_csr_translator:uav_lock
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_read -> sgdma_tx_csr_translator:uav_read
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0);  -- sgdma_tx_csr_translator:uav_readdata -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                      -- sgdma_tx_csr_translator:uav_readdatavalid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sgdma_tx_csr_translator:uav_debugaccess
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);   -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> sgdma_tx_csr_translator:uav_byteenable
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(94 downto 0);  -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(94 downto 0);  -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0);  -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                      -- sgdma_rx_csr_translator:uav_waitrequest -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);   -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_burstcount -> sgdma_rx_csr_translator:uav_burstcount
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0);  -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_writedata -> sgdma_rx_csr_translator:uav_writedata
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(22 downto 0);  -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_address -> sgdma_rx_csr_translator:uav_address
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_write -> sgdma_rx_csr_translator:uav_write
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_lock -> sgdma_rx_csr_translator:uav_lock
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_read -> sgdma_rx_csr_translator:uav_read
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0);  -- sgdma_rx_csr_translator:uav_readdata -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                      -- sgdma_rx_csr_translator:uav_readdatavalid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sgdma_rx_csr_translator:uav_debugaccess
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);   -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:m0_byteenable -> sgdma_rx_csr_translator:uav_byteenable
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(94 downto 0);  -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(94 downto 0);  -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0);  -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_waitrequest                                  : std_logic;                      -- cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_to_flash_ccb_m0_translator:uav_waitrequest
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_burstcount                                   : std_logic_vector(2 downto 0);   -- cpu_to_flash_ccb_m0_translator:uav_burstcount -> cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_writedata                                    : std_logic_vector(31 downto 0);  -- cpu_to_flash_ccb_m0_translator:uav_writedata -> cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_address                                      : std_logic_vector(27 downto 0);  -- cpu_to_flash_ccb_m0_translator:uav_address -> cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:av_address
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_lock                                         : std_logic;                      -- cpu_to_flash_ccb_m0_translator:uav_lock -> cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_write                                        : std_logic;                      -- cpu_to_flash_ccb_m0_translator:uav_write -> cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:av_write
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_read                                         : std_logic;                      -- cpu_to_flash_ccb_m0_translator:uav_read -> cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:av_read
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_readdata                                     : std_logic_vector(31 downto 0);  -- cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:av_readdata -> cpu_to_flash_ccb_m0_translator:uav_readdata
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_debugaccess                                  : std_logic;                      -- cpu_to_flash_ccb_m0_translator:uav_debugaccess -> cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_byteenable                                   : std_logic_vector(3 downto 0);   -- cpu_to_flash_ccb_m0_translator:uav_byteenable -> cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_readdatavalid                                : std_logic;                      -- cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_to_flash_ccb_m0_translator:uav_readdatavalid
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator:uav_waitrequest -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(1 downto 0);   -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> cfi_flash_ts_controller_fpga_uas_translator:uav_burstcount
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(15 downto 0);  -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> cfi_flash_ts_controller_fpga_uas_translator:uav_writedata
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(27 downto 0);  -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:m0_address -> cfi_flash_ts_controller_fpga_uas_translator:uav_address
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:m0_write -> cfi_flash_ts_controller_fpga_uas_translator:uav_write
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:m0_lock -> cfi_flash_ts_controller_fpga_uas_translator:uav_lock
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:m0_read -> cfi_flash_ts_controller_fpga_uas_translator:uav_read
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(15 downto 0);  -- cfi_flash_ts_controller_fpga_uas_translator:uav_readdata -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator:uav_readdatavalid -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cfi_flash_ts_controller_fpga_uas_translator:uav_debugaccess
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(1 downto 0);   -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> cfi_flash_ts_controller_fpga_uas_translator:uav_byteenable
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(77 downto 0);  -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(77 downto 0);  -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(17 downto 0);  -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid       : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data        : std_logic_vector(17 downto 0);  -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready       : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest                  : std_logic;                      -- cfi_flash_ts_controller_uas_translator:uav_waitrequest -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_burstcount                   : std_logic_vector(1 downto 0);   -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> cfi_flash_ts_controller_uas_translator:uav_burstcount
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_writedata                    : std_logic_vector(15 downto 0);  -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> cfi_flash_ts_controller_uas_translator:uav_writedata
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_address                      : std_logic_vector(27 downto 0);  -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:m0_address -> cfi_flash_ts_controller_uas_translator:uav_address
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_write                        : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:m0_write -> cfi_flash_ts_controller_uas_translator:uav_write
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_lock                         : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:m0_lock -> cfi_flash_ts_controller_uas_translator:uav_lock
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_read                         : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:m0_read -> cfi_flash_ts_controller_uas_translator:uav_read
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_readdata                     : std_logic_vector(15 downto 0);  -- cfi_flash_ts_controller_uas_translator:uav_readdata -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid                : std_logic;                      -- cfi_flash_ts_controller_uas_translator:uav_readdatavalid -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess                  : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cfi_flash_ts_controller_uas_translator:uav_debugaccess
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_byteenable                   : std_logic_vector(1 downto 0);   -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> cfi_flash_ts_controller_uas_translator:uav_byteenable
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket           : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_valid                 : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket         : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_data                  : std_logic_vector(77 downto 0);  -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_ready                 : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket        : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid              : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket      : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data               : std_logic_vector(77 downto 0);  -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready              : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid            : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data             : std_logic_vector(17 downto 0);  -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready            : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid            : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data             : std_logic_vector(17 downto 0);  -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready            : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest                                      : std_logic;                      -- sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_tx_m_read_translator:uav_waitrequest
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount                                       : std_logic_vector(2 downto 0);   -- sgdma_tx_m_read_translator:uav_burstcount -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_burstcount
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_writedata                                        : std_logic_vector(31 downto 0);  -- sgdma_tx_m_read_translator:uav_writedata -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_writedata
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_address                                          : std_logic_vector(31 downto 0);  -- sgdma_tx_m_read_translator:uav_address -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_address
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_lock                                             : std_logic;                      -- sgdma_tx_m_read_translator:uav_lock -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_lock
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_write                                            : std_logic;                      -- sgdma_tx_m_read_translator:uav_write -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_write
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_read                                             : std_logic;                      -- sgdma_tx_m_read_translator:uav_read -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_read
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_readdata                                         : std_logic_vector(31 downto 0);  -- sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_tx_m_read_translator:uav_readdata
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess                                      : std_logic;                      -- sgdma_tx_m_read_translator:uav_debugaccess -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_debugaccess
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable                                       : std_logic_vector(3 downto 0);   -- sgdma_tx_m_read_translator:uav_byteenable -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_byteenable
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid                                    : std_logic;                      -- sgdma_tx_m_read_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_tx_m_read_translator:uav_readdatavalid
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest                                     : std_logic;                      -- sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_waitrequest -> sgdma_rx_m_write_translator:uav_waitrequest
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount                                      : std_logic_vector(2 downto 0);   -- sgdma_rx_m_write_translator:uav_burstcount -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_burstcount
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_writedata                                       : std_logic_vector(31 downto 0);  -- sgdma_rx_m_write_translator:uav_writedata -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_writedata
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_address                                         : std_logic_vector(31 downto 0);  -- sgdma_rx_m_write_translator:uav_address -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_address
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_lock                                            : std_logic;                      -- sgdma_rx_m_write_translator:uav_lock -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_lock
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_write                                           : std_logic;                      -- sgdma_rx_m_write_translator:uav_write -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_write
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_read                                            : std_logic;                      -- sgdma_rx_m_write_translator:uav_read -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_read
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_readdata                                        : std_logic_vector(31 downto 0);  -- sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_readdata -> sgdma_rx_m_write_translator:uav_readdata
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess                                     : std_logic;                      -- sgdma_rx_m_write_translator:uav_debugaccess -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_debugaccess
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable                                      : std_logic_vector(3 downto 0);   -- sgdma_rx_m_write_translator:uav_byteenable -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_byteenable
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid                                   : std_logic;                      -- sgdma_rx_m_write_translator_avalon_universal_master_0_agent:av_readdatavalid -> sgdma_rx_m_write_translator:uav_readdatavalid
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest                      : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator:uav_waitrequest -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount                       : std_logic_vector(2 downto 0);   -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> tse_dma_to_sdram_ccb_s0_translator:uav_burstcount
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_writedata                        : std_logic_vector(31 downto 0);  -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> tse_dma_to_sdram_ccb_s0_translator:uav_writedata
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_address                          : std_logic_vector(31 downto 0);  -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:m0_address -> tse_dma_to_sdram_ccb_s0_translator:uav_address
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_write                            : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:m0_write -> tse_dma_to_sdram_ccb_s0_translator:uav_write
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_lock                             : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:m0_lock -> tse_dma_to_sdram_ccb_s0_translator:uav_lock
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_read                             : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:m0_read -> tse_dma_to_sdram_ccb_s0_translator:uav_read
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdata                         : std_logic_vector(31 downto 0);  -- tse_dma_to_sdram_ccb_s0_translator:uav_readdata -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                    : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator:uav_readdatavalid -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess                      : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> tse_dma_to_sdram_ccb_s0_translator:uav_debugaccess
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable                       : std_logic_vector(3 downto 0);   -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> tse_dma_to_sdram_ccb_s0_translator:uav_byteenable
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket               : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid                     : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket             : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_data                      : std_logic_vector(99 downto 0);  -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready                     : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket            : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                  : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket          : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                   : std_logic_vector(99 downto 0);  -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                  : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                 : std_logic_vector(33 downto 0);  -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_waitrequest                              : std_logic;                      -- tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> tse_dma_to_sdram_ccb_m0_translator:uav_waitrequest
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_burstcount                               : std_logic_vector(2 downto 0);   -- tse_dma_to_sdram_ccb_m0_translator:uav_burstcount -> tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:av_burstcount
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_writedata                                : std_logic_vector(31 downto 0);  -- tse_dma_to_sdram_ccb_m0_translator:uav_writedata -> tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:av_writedata
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_address                                  : std_logic_vector(26 downto 0);  -- tse_dma_to_sdram_ccb_m0_translator:uav_address -> tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:av_address
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_lock                                     : std_logic;                      -- tse_dma_to_sdram_ccb_m0_translator:uav_lock -> tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:av_lock
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_write                                    : std_logic;                      -- tse_dma_to_sdram_ccb_m0_translator:uav_write -> tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:av_write
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_read                                     : std_logic;                      -- tse_dma_to_sdram_ccb_m0_translator:uav_read -> tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:av_read
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_readdata                                 : std_logic_vector(31 downto 0);  -- tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:av_readdata -> tse_dma_to_sdram_ccb_m0_translator:uav_readdata
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_debugaccess                              : std_logic;                      -- tse_dma_to_sdram_ccb_m0_translator:uav_debugaccess -> tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_byteenable                               : std_logic_vector(3 downto 0);   -- tse_dma_to_sdram_ccb_m0_translator:uav_byteenable -> tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:av_byteenable
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_readdatavalid                            : std_logic;                      -- tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> tse_dma_to_sdram_ccb_m0_translator:uav_readdatavalid
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_waitrequest                                   : std_logic;                      -- cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_to_sdram_pb_m0_translator:uav_waitrequest
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_burstcount                                    : std_logic_vector(2 downto 0);   -- cpu_to_sdram_pb_m0_translator:uav_burstcount -> cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_writedata                                     : std_logic_vector(31 downto 0);  -- cpu_to_sdram_pb_m0_translator:uav_writedata -> cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_address                                       : std_logic_vector(26 downto 0);  -- cpu_to_sdram_pb_m0_translator:uav_address -> cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:av_address
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_lock                                          : std_logic;                      -- cpu_to_sdram_pb_m0_translator:uav_lock -> cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_write                                         : std_logic;                      -- cpu_to_sdram_pb_m0_translator:uav_write -> cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:av_write
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_read                                          : std_logic;                      -- cpu_to_sdram_pb_m0_translator:uav_read -> cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:av_read
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_readdata                                      : std_logic_vector(31 downto 0);  -- cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:av_readdata -> cpu_to_sdram_pb_m0_translator:uav_readdata
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_debugaccess                                   : std_logic;                      -- cpu_to_sdram_pb_m0_translator:uav_debugaccess -> cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_byteenable                                    : std_logic_vector(3 downto 0);   -- cpu_to_sdram_pb_m0_translator:uav_byteenable -> cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_readdatavalid                                 : std_logic;                      -- cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_to_sdram_pb_m0_translator:uav_readdatavalid
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest                                  : std_logic;                      -- sdram_0_avl_translator:uav_waitrequest -> sdram_0_avl_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_burstcount                                   : std_logic_vector(5 downto 0);   -- sdram_0_avl_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_0_avl_translator:uav_burstcount
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_writedata                                    : std_logic_vector(63 downto 0);  -- sdram_0_avl_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_0_avl_translator:uav_writedata
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_address                                      : std_logic_vector(26 downto 0);  -- sdram_0_avl_translator_avalon_universal_slave_0_agent:m0_address -> sdram_0_avl_translator:uav_address
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_write                                        : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent:m0_write -> sdram_0_avl_translator:uav_write
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_lock                                         : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_0_avl_translator:uav_lock
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_read                                         : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent:m0_read -> sdram_0_avl_translator:uav_read
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_readdata                                     : std_logic_vector(63 downto 0);  -- sdram_0_avl_translator:uav_readdata -> sdram_0_avl_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                : std_logic;                      -- sdram_0_avl_translator:uav_readdatavalid -> sdram_0_avl_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess                                  : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_0_avl_translator:uav_debugaccess
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_byteenable                                   : std_logic_vector(7 downto 0);   -- sdram_0_avl_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_0_avl_translator:uav_byteenable
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                           : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rf_source_valid                                 : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                         : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rf_source_data                                  : std_logic_vector(133 downto 0); -- sdram_0_avl_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rf_source_ready                                 : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_0_avl_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                        : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                              : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                      : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                               : std_logic_vector(133 downto 0); -- sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                              : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                            : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                             : std_logic_vector(65 downto 0);  -- sdram_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                            : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_0_avl_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal linux_cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                       : std_logic;                      -- linux_cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal linux_cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid                             : std_logic;                      -- linux_cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal linux_cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                     : std_logic;                      -- linux_cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal linux_cpu_data_master_translator_avalon_universal_master_0_agent_cp_data                              : std_logic_vector(99 downto 0);  -- linux_cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal linux_cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready                             : std_logic;                      -- addr_router:sink_ready -> linux_cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket                : std_logic;                      -- linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                      : std_logic;                      -- linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket              : std_logic;                      -- linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data                       : std_logic_vector(99 downto 0);  -- linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal linux_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                      : std_logic;                      -- addr_router_001:sink_ready -> linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket                  : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                        : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket                : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                         : std_logic_vector(99 downto 0);  -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                        : std_logic;                      -- id_router:sink_ready -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket                          : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rp_valid                                : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket                        : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rp_data                                 : std_logic_vector(99 downto 0);  -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rp_ready                                : std_logic;                      -- id_router_001:sink_ready -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:rp_ready
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket                    : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rp_valid                          : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket                  : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rp_data                           : std_logic_vector(99 downto 0);  -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rp_ready                          : std_logic;                      -- id_router_002:sink_ready -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:rp_ready
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket                           : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rp_valid                                 : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket                         : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rp_data                                  : std_logic_vector(99 downto 0);  -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rp_ready                                 : std_logic;                      -- id_router_003:sink_ready -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:rp_ready
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket                   : std_logic;                      -- sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid                         : std_logic;                      -- sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket                 : std_logic;                      -- sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data                          : std_logic_vector(100 downto 0); -- sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	signal sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready                         : std_logic;                      -- addr_router_002:sink_ready -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:cp_ready
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket                   : std_logic;                      -- sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid                         : std_logic;                      -- sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket                 : std_logic;                      -- sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data                          : std_logic_vector(100 downto 0); -- sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	signal sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready                         : std_logic;                      -- addr_router_003:sink_ready -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:cp_ready
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket                    : std_logic;                      -- sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid                          : std_logic;                      -- sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket                  : std_logic;                      -- sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data                           : std_logic_vector(100 downto 0); -- sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	signal sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready                          : std_logic;                      -- addr_router_004:sink_ready -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:cp_ready
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket                    : std_logic;                      -- sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid                          : std_logic;                      -- sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket                  : std_logic;                      -- sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data                           : std_logic_vector(100 downto 0); -- sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	signal sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready                          : std_logic;                      -- addr_router_005:sink_ready -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:cp_ready
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket                     : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rp_valid                           : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket                   : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rp_data                            : std_logic_vector(100 downto 0); -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rp_ready                           : std_logic;                      -- id_router_004:sink_ready -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:rp_ready
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent_cp_endofpacket                    : std_logic;                      -- dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_006:sink_endofpacket
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent_cp_valid                          : std_logic;                      -- dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_006:sink_valid
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent_cp_startofpacket                  : std_logic;                      -- dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_006:sink_startofpacket
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent_cp_data                           : std_logic_vector(93 downto 0);  -- dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_006:sink_data
	signal dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent_cp_ready                          : std_logic;                      -- addr_router_006:sink_ready -> dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket                   : std_logic;                      -- cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_007:sink_endofpacket
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent_cp_valid                         : std_logic;                      -- cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_007:sink_valid
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket                 : std_logic;                      -- cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_007:sink_startofpacket
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent_cp_data                          : std_logic_vector(93 downto 0);  -- cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_007:sink_data
	signal cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent_cp_ready                         : std_logic;                      -- addr_router_007:sink_ready -> cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:cp_ready
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                         : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid                               : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                       : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data                                : std_logic_vector(93 downto 0);  -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready                               : std_logic;                      -- id_router_005:sink_ready -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                  : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                        : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                         : std_logic_vector(93 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                        : std_logic;                      -- id_router_006:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket                         : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid                               : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket                       : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data                                : std_logic_vector(93 downto 0);  -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready                               : std_logic;                      -- id_router_007:sink_ready -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                          : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                                : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                        : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data                                 : std_logic_vector(93 downto 0);  -- sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	signal sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                                : std_logic;                      -- id_router_008:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                           : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rp_valid                                 : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                         : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rp_data                                  : std_logic_vector(93 downto 0);  -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	signal linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rp_ready                                 : std_logic;                      -- id_router_009:sink_ready -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket                               : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rp_valid                                     : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket                             : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rp_data                                      : std_logic_vector(93 downto 0);  -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	signal gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rp_ready                                     : std_logic;                      -- id_router_010:sink_ready -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:rp_ready
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(93 downto 0);  -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	signal sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                      -- id_router_011:sink_ready -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:rp_ready
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(93 downto 0);  -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	signal sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                      -- id_router_012:sink_ready -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:rp_ready
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket                         : std_logic;                      -- cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_008:sink_endofpacket
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent_cp_valid                               : std_logic;                      -- cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_008:sink_valid
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket                       : std_logic;                      -- cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_008:sink_startofpacket
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent_cp_data                                : std_logic_vector(94 downto 0);  -- cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_008:sink_data
	signal cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent_cp_ready                               : std_logic;                      -- addr_router_008:sink_ready -> cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:cp_ready
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(76 downto 0);  -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	signal cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                      -- id_router_013:sink_ready -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:rp_ready
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket                  : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rp_valid                        : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket                : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rp_data                         : std_logic_vector(76 downto 0);  -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	signal cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rp_ready                        : std_logic;                      -- id_router_014:sink_ready -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:rp_ready
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket                             : std_logic;                      -- sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_009:sink_endofpacket
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid                                   : std_logic;                      -- sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_009:sink_valid
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket                           : std_logic;                      -- sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_009:sink_startofpacket
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data                                    : std_logic_vector(98 downto 0);  -- sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_data -> addr_router_009:sink_data
	signal sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready                                   : std_logic;                      -- addr_router_009:sink_ready -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:cp_ready
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket                            : std_logic;                      -- sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_010:sink_endofpacket
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid                                  : std_logic;                      -- sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_010:sink_valid
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket                          : std_logic;                      -- sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_010:sink_startofpacket
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data                                   : std_logic_vector(98 downto 0);  -- sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_data -> addr_router_010:sink_data
	signal sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready                                  : std_logic;                      -- addr_router_010:sink_ready -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:cp_ready
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket                      : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rp_valid                            : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket                    : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rp_data                             : std_logic_vector(98 downto 0);  -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	signal tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rp_ready                            : std_logic;                      -- id_router_015:sink_ready -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:rp_ready
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket                     : std_logic;                      -- tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_011:sink_endofpacket
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent_cp_valid                           : std_logic;                      -- tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_011:sink_valid
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket                   : std_logic;                      -- tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_011:sink_startofpacket
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent_cp_data                            : std_logic_vector(96 downto 0);  -- tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_011:sink_data
	signal tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent_cp_ready                           : std_logic;                      -- addr_router_011:sink_ready -> tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket                          : std_logic;                      -- cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_012:sink_endofpacket
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent_cp_valid                                : std_logic;                      -- cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_012:sink_valid
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket                        : std_logic;                      -- cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_012:sink_startofpacket
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent_cp_data                                 : std_logic_vector(96 downto 0);  -- cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_012:sink_data
	signal cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent_cp_ready                                : std_logic;                      -- addr_router_012:sink_ready -> cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:cp_ready
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket                                  : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rp_valid                                        : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket                                : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rp_data                                         : std_logic_vector(132 downto 0); -- sdram_0_avl_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	signal sdram_0_avl_translator_avalon_universal_slave_0_agent_rp_ready                                        : std_logic;                      -- id_router_016:sink_ready -> sdram_0_avl_translator_avalon_universal_slave_0_agent:rp_ready
	signal addr_router_src_endofpacket                                                                           : std_logic;                      -- addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	signal addr_router_src_valid                                                                                 : std_logic;                      -- addr_router:src_valid -> limiter:cmd_sink_valid
	signal addr_router_src_startofpacket                                                                         : std_logic;                      -- addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	signal addr_router_src_data                                                                                  : std_logic_vector(99 downto 0);  -- addr_router:src_data -> limiter:cmd_sink_data
	signal addr_router_src_channel                                                                               : std_logic_vector(3 downto 0);   -- addr_router:src_channel -> limiter:cmd_sink_channel
	signal addr_router_src_ready                                                                                 : std_logic;                      -- limiter:cmd_sink_ready -> addr_router:src_ready
	signal limiter_rsp_src_endofpacket                                                                           : std_logic;                      -- limiter:rsp_src_endofpacket -> linux_cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_rsp_src_valid                                                                                 : std_logic;                      -- limiter:rsp_src_valid -> linux_cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_rsp_src_startofpacket                                                                         : std_logic;                      -- limiter:rsp_src_startofpacket -> linux_cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_rsp_src_data                                                                                  : std_logic_vector(99 downto 0);  -- limiter:rsp_src_data -> linux_cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_rsp_src_channel                                                                               : std_logic_vector(3 downto 0);   -- limiter:rsp_src_channel -> linux_cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_rsp_src_ready                                                                                 : std_logic;                      -- linux_cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	signal addr_router_001_src_endofpacket                                                                       : std_logic;                      -- addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	signal addr_router_001_src_valid                                                                             : std_logic;                      -- addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	signal addr_router_001_src_startofpacket                                                                     : std_logic;                      -- addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	signal addr_router_001_src_data                                                                              : std_logic_vector(99 downto 0);  -- addr_router_001:src_data -> limiter_001:cmd_sink_data
	signal addr_router_001_src_channel                                                                           : std_logic_vector(3 downto 0);   -- addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	signal addr_router_001_src_ready                                                                             : std_logic;                      -- limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	signal limiter_001_rsp_src_endofpacket                                                                       : std_logic;                      -- limiter_001:rsp_src_endofpacket -> linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_001_rsp_src_valid                                                                             : std_logic;                      -- limiter_001:rsp_src_valid -> linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_001_rsp_src_startofpacket                                                                     : std_logic;                      -- limiter_001:rsp_src_startofpacket -> linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_001_rsp_src_data                                                                              : std_logic_vector(99 downto 0);  -- limiter_001:rsp_src_data -> linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_001_rsp_src_channel                                                                           : std_logic_vector(3 downto 0);   -- limiter_001:rsp_src_channel -> linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_001_rsp_src_ready                                                                             : std_logic;                      -- linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	signal addr_router_007_src_endofpacket                                                                       : std_logic;                      -- addr_router_007:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	signal addr_router_007_src_valid                                                                             : std_logic;                      -- addr_router_007:src_valid -> limiter_002:cmd_sink_valid
	signal addr_router_007_src_startofpacket                                                                     : std_logic;                      -- addr_router_007:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	signal addr_router_007_src_data                                                                              : std_logic_vector(93 downto 0);  -- addr_router_007:src_data -> limiter_002:cmd_sink_data
	signal addr_router_007_src_channel                                                                           : std_logic_vector(7 downto 0);   -- addr_router_007:src_channel -> limiter_002:cmd_sink_channel
	signal addr_router_007_src_ready                                                                             : std_logic;                      -- limiter_002:cmd_sink_ready -> addr_router_007:src_ready
	signal limiter_002_rsp_src_endofpacket                                                                       : std_logic;                      -- limiter_002:rsp_src_endofpacket -> cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_002_rsp_src_valid                                                                             : std_logic;                      -- limiter_002:rsp_src_valid -> cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_002_rsp_src_startofpacket                                                                     : std_logic;                      -- limiter_002:rsp_src_startofpacket -> cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_002_rsp_src_data                                                                              : std_logic_vector(93 downto 0);  -- limiter_002:rsp_src_data -> cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_002_rsp_src_channel                                                                           : std_logic_vector(7 downto 0);   -- limiter_002:rsp_src_channel -> cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_002_rsp_src_ready                                                                             : std_logic;                      -- cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_002:rsp_src_ready
	signal addr_router_008_src_endofpacket                                                                       : std_logic;                      -- addr_router_008:src_endofpacket -> limiter_003:cmd_sink_endofpacket
	signal addr_router_008_src_valid                                                                             : std_logic;                      -- addr_router_008:src_valid -> limiter_003:cmd_sink_valid
	signal addr_router_008_src_startofpacket                                                                     : std_logic;                      -- addr_router_008:src_startofpacket -> limiter_003:cmd_sink_startofpacket
	signal addr_router_008_src_data                                                                              : std_logic_vector(94 downto 0);  -- addr_router_008:src_data -> limiter_003:cmd_sink_data
	signal addr_router_008_src_channel                                                                           : std_logic_vector(1 downto 0);   -- addr_router_008:src_channel -> limiter_003:cmd_sink_channel
	signal addr_router_008_src_ready                                                                             : std_logic;                      -- limiter_003:cmd_sink_ready -> addr_router_008:src_ready
	signal limiter_003_rsp_src_endofpacket                                                                       : std_logic;                      -- limiter_003:rsp_src_endofpacket -> cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_003_rsp_src_valid                                                                             : std_logic;                      -- limiter_003:rsp_src_valid -> cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_003_rsp_src_startofpacket                                                                     : std_logic;                      -- limiter_003:rsp_src_startofpacket -> cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_003_rsp_src_data                                                                              : std_logic_vector(94 downto 0);  -- limiter_003:rsp_src_data -> cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_003_rsp_src_channel                                                                           : std_logic_vector(1 downto 0);   -- limiter_003:rsp_src_channel -> cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_003_rsp_src_ready                                                                             : std_logic;                      -- cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_003:rsp_src_ready
	signal burst_adapter_source0_endofpacket                                                                     : std_logic;                      -- burst_adapter:source0_endofpacket -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_source0_valid                                                                           : std_logic;                      -- burst_adapter:source0_valid -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_source0_startofpacket                                                                   : std_logic;                      -- burst_adapter:source0_startofpacket -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_source0_data                                                                            : std_logic_vector(76 downto 0);  -- burst_adapter:source0_data -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_source0_ready                                                                           : std_logic;                      -- cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	signal burst_adapter_source0_channel                                                                         : std_logic_vector(1 downto 0);   -- burst_adapter:source0_channel -> cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_001_source0_endofpacket                                                                 : std_logic;                      -- burst_adapter_001:source0_endofpacket -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_001_source0_valid                                                                       : std_logic;                      -- burst_adapter_001:source0_valid -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_001_source0_startofpacket                                                               : std_logic;                      -- burst_adapter_001:source0_startofpacket -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_001_source0_data                                                                        : std_logic_vector(76 downto 0);  -- burst_adapter_001:source0_data -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_001_source0_ready                                                                       : std_logic;                      -- cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	signal burst_adapter_001_source0_channel                                                                     : std_logic_vector(1 downto 0);   -- burst_adapter_001:source0_channel -> cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:cp_channel
	signal rst_controller_reset_out_reset                                                                        : std_logic;                      -- rst_controller:reset_out -> [addr_router_002:reset, addr_router_003:reset, addr_router_004:reset, addr_router_005:reset, addr_router_006:reset, addr_router_007:reset, addr_router_008:reset, addr_router_009:reset, addr_router_010:reset, avalon_st_adapter:in_rst_0_reset, burst_adapter:reset, burst_adapter_001:reset, cfi_flash_ts_bridge:reset, cfi_flash_ts_bridge_fpga:reset, cfi_flash_ts_controller:reset_reset, cfi_flash_ts_controller_fpga:reset_reset, cfi_flash_ts_controller_fpga_uas_translator:reset, cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent:reset, cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cfi_flash_ts_controller_uas_translator:reset, cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent:reset, cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux_002:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_demux_005:reset, cmd_xbar_demux_006:reset, cmd_xbar_demux_007:reset, cmd_xbar_demux_008:reset, cmd_xbar_demux_009:reset, cmd_xbar_demux_010:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_015:reset, cpu_to_flash_ccb:m0_reset, cpu_to_flash_ccb_m0_translator:reset, cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent:reset, cpu_to_peripherals_ccb:m0_reset, cpu_to_peripherals_ccb_m0_translator:reset, cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent:reset, descriptor_memory:reset, descriptor_memory_s1_translator:reset, descriptor_memory_s1_translator_avalon_universal_slave_0_agent:reset, descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dma_to_descriptor_mem:reset, dma_to_descriptor_mem_m0_translator:reset, dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:reset, dma_to_descriptor_mem_s0_translator:reset, dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:reset, dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, gtp_regif_0_s0_translator:reset, gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:reset, gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter_002:reset, limiter_003:reset, linux_timer_1ms_s1_translator:reset, linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:reset, linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_mux_007:reset, rsp_xbar_mux_008:reset, rst_controller_reset_out_reset:in, sgdma_rx_csr_translator:reset, sgdma_rx_csr_translator_avalon_universal_slave_0_agent:reset, sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_rx_descriptor_read_translator:reset, sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:reset, sgdma_rx_descriptor_write_translator:reset, sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:reset, sgdma_rx_m_write_translator:reset, sgdma_rx_m_write_translator_avalon_universal_master_0_agent:reset, sgdma_tx_csr_translator:reset, sgdma_tx_csr_translator_avalon_universal_slave_0_agent:reset, sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sgdma_tx_descriptor_read_translator:reset, sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:reset, sgdma_tx_descriptor_write_translator:reset, sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:reset, sgdma_tx_m_read_translator:reset, sgdma_tx_m_read_translator_avalon_universal_master_0_agent:reset, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, tse_dma_to_sdram_ccb:s0_reset, tse_dma_to_sdram_ccb_s0_translator:reset, tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:reset, tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, tse_mac:reset, tse_mac_control_port_translator:reset, tse_mac_control_port_translator_avalon_universal_slave_0_agent:reset, tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset]
	signal rst_controller_reset_out_reset_req                                                                    : std_logic;                      -- rst_controller:reset_req -> descriptor_memory:reset_req
	signal linux_cpu_jtag_debug_module_reset_reset                                                               : std_logic;                      -- linux_cpu:jtag_debug_module_resetrequest -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in1, rst_controller_003:reset_in2]
	signal sdram_0_afi_reset_reset                                                                               : std_logic;                      -- sdram_0:afi_reset_n -> sdram_0_afi_reset_reset:in
	signal rst_controller_001_reset_out_reset                                                                    : std_logic;                      -- rst_controller_001:reset_out -> [addr_router:reset, addr_router_001:reset, addr_router_011:reset, addr_router_012:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_011:reset, cmd_xbar_demux_012:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_003:reset, cpu_to_flash_ccb:s0_reset, cpu_to_flash_ccb_s0_translator:reset, cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:reset, cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cpu_to_peripherals_ccb:s0_reset, cpu_to_peripherals_ccb_s0_translator:reset, cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:reset, cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cpu_to_sdram_pb:reset, cpu_to_sdram_pb_m0_translator:reset, cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:reset, cpu_to_sdram_pb_s0_translator:reset, cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:reset, cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, limiter:reset, limiter_001:reset, linux_cpu_data_master_translator:reset, linux_cpu_data_master_translator_avalon_universal_master_0_agent:reset, linux_cpu_instruction_master_translator:reset, linux_cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, linux_cpu_jtag_debug_module_translator:reset, linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, linux_cpu_tightly_coupled_data_master_0_translator:reset, linux_cpu_tightly_coupled_instruction_master_0_translator:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_001_reset_out_reset:in, tlb_miss_ram_1k:reset, tlb_miss_ram_1k:reset2, tlb_miss_ram_1k_s1_translator:reset, tlb_miss_ram_1k_s2_translator:reset, tse_dma_to_sdram_ccb:m0_reset, tse_dma_to_sdram_ccb_m0_translator:reset, tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:reset]
	signal rst_controller_001_reset_out_reset_req                                                                : std_logic;                      -- rst_controller_001:reset_req -> [tlb_miss_ram_1k:reset_req, tlb_miss_ram_1k:reset_req2]
	signal rst_controller_002_reset_out_reset                                                                    : std_logic;                      -- rst_controller_002:reset_out -> rst_controller_002_reset_out_reset:in
	signal rst_controller_003_reset_out_reset                                                                    : std_logic;                      -- rst_controller_003:reset_out -> [gtp_regif_0:reset, irq_synchronizer_004:receiver_reset]
	signal rst_controller_004_reset_out_reset                                                                    : std_logic;                      -- rst_controller_004:reset_out -> [cmd_xbar_mux_016:reset, id_router_016:reset, rsp_xbar_demux_016:reset, sdram_0_avl_translator:reset, sdram_0_avl_translator_avalon_universal_slave_0_agent:reset, sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter_004:reset, width_adapter_005:reset]
	signal cmd_xbar_demux_src0_endofpacket                                                                       : std_logic;                      -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                             : std_logic;                      -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                           : std_logic_vector(3 downto 0);   -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                             : std_logic;                      -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                       : std_logic;                      -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                             : std_logic;                      -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                           : std_logic_vector(3 downto 0);   -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                             : std_logic;                      -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_src2_endofpacket                                                                       : std_logic;                      -- cmd_xbar_demux:src2_endofpacket -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_src2_valid                                                                             : std_logic;                      -- cmd_xbar_demux:src2_valid -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_src2_startofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src2_startofpacket -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_src2_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src2_data -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_src2_channel                                                                           : std_logic_vector(3 downto 0);   -- cmd_xbar_demux:src2_channel -> cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_src3_endofpacket                                                                       : std_logic;                      -- cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	signal cmd_xbar_demux_src3_valid                                                                             : std_logic;                      -- cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	signal cmd_xbar_demux_src3_startofpacket                                                                     : std_logic;                      -- cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	signal cmd_xbar_demux_src3_data                                                                              : std_logic_vector(99 downto 0);  -- cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	signal cmd_xbar_demux_src3_channel                                                                           : std_logic_vector(3 downto 0);   -- cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	signal cmd_xbar_demux_src3_ready                                                                             : std_logic;                      -- cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                          : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                       : std_logic_vector(3 downto 0);   -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                         : std_logic;                      -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                          : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                       : std_logic_vector(3 downto 0);   -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                         : std_logic;                      -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src2_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_003:sink1_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                          : std_logic_vector(99 downto 0);  -- cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_003:sink1_data
	signal cmd_xbar_demux_001_src2_channel                                                                       : std_logic_vector(3 downto 0);   -- cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_003:sink1_channel
	signal cmd_xbar_demux_001_src2_ready                                                                         : std_logic;                      -- cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src2_ready
	signal rsp_xbar_demux_src0_endofpacket                                                                       : std_logic;                      -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                             : std_logic;                      -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                     : std_logic;                      -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                              : std_logic_vector(99 downto 0);  -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                           : std_logic_vector(3 downto 0);   -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                             : std_logic;                      -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                       : std_logic;                      -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                             : std_logic;                      -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                     : std_logic;                      -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                              : std_logic_vector(99 downto 0);  -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                           : std_logic_vector(3 downto 0);   -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                             : std_logic;                      -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                          : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                       : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                         : std_logic;                      -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                         : std_logic;                      -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                          : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                                       : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                         : std_logic;                      -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                          : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                                       : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                         : std_logic;                      -- rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                          : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	signal rsp_xbar_demux_003_src0_channel                                                                       : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	signal rsp_xbar_demux_003_src0_ready                                                                         : std_logic;                      -- rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	signal rsp_xbar_demux_003_src1_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal rsp_xbar_demux_003_src1_valid                                                                         : std_logic;                      -- rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink2_valid
	signal rsp_xbar_demux_003_src1_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal rsp_xbar_demux_003_src1_data                                                                          : std_logic_vector(99 downto 0);  -- rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink2_data
	signal rsp_xbar_demux_003_src1_channel                                                                       : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_003_src1_ready                                                                         : std_logic;                      -- rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_003:src1_ready
	signal limiter_cmd_src_endofpacket                                                                           : std_logic;                      -- limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal limiter_cmd_src_startofpacket                                                                         : std_logic;                      -- limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal limiter_cmd_src_data                                                                                  : std_logic_vector(99 downto 0);  -- limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	signal limiter_cmd_src_channel                                                                               : std_logic_vector(3 downto 0);   -- limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	signal limiter_cmd_src_ready                                                                                 : std_logic;                      -- cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                          : std_logic;                      -- rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	signal rsp_xbar_mux_src_valid                                                                                : std_logic;                      -- rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	signal rsp_xbar_mux_src_startofpacket                                                                        : std_logic;                      -- rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	signal rsp_xbar_mux_src_data                                                                                 : std_logic_vector(99 downto 0);  -- rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	signal rsp_xbar_mux_src_channel                                                                              : std_logic_vector(3 downto 0);   -- rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	signal rsp_xbar_mux_src_ready                                                                                : std_logic;                      -- limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	signal limiter_001_cmd_src_endofpacket                                                                       : std_logic;                      -- limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal limiter_001_cmd_src_startofpacket                                                                     : std_logic;                      -- limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal limiter_001_cmd_src_data                                                                              : std_logic_vector(99 downto 0);  -- limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	signal limiter_001_cmd_src_channel                                                                           : std_logic_vector(3 downto 0);   -- limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	signal limiter_001_cmd_src_ready                                                                             : std_logic;                      -- cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                      : std_logic;                      -- rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                            : std_logic;                      -- rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                                    : std_logic;                      -- rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                             : std_logic_vector(99 downto 0);  -- rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	signal rsp_xbar_mux_001_src_channel                                                                          : std_logic_vector(3 downto 0);   -- rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	signal rsp_xbar_mux_001_src_ready                                                                            : std_logic;                      -- limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	signal cmd_xbar_mux_src_endofpacket                                                                          : std_logic;                      -- cmd_xbar_mux:src_endofpacket -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_src_valid                                                                                : std_logic;                      -- cmd_xbar_mux:src_valid -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_src_startofpacket                                                                        : std_logic;                      -- cmd_xbar_mux:src_startofpacket -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_src_data                                                                                 : std_logic_vector(99 downto 0);  -- cmd_xbar_mux:src_data -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_src_channel                                                                              : std_logic_vector(3 downto 0);   -- cmd_xbar_mux:src_channel -> linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_src_ready                                                                                : std_logic;                      -- linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                             : std_logic;                      -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                                   : std_logic;                      -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                           : std_logic;                      -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                                    : std_logic_vector(99 downto 0);  -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                                 : std_logic_vector(3 downto 0);   -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                                   : std_logic;                      -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                      : std_logic;                      -- cmd_xbar_mux_001:src_endofpacket -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                            : std_logic;                      -- cmd_xbar_mux_001:src_valid -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_001:src_startofpacket -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                             : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_001:src_data -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_001_src_channel                                                                          : std_logic_vector(3 downto 0);   -- cmd_xbar_mux_001:src_channel -> cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_001_src_ready                                                                            : std_logic;                      -- cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	signal id_router_001_src_endofpacket                                                                         : std_logic;                      -- id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal id_router_001_src_valid                                                                               : std_logic;                      -- id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	signal id_router_001_src_startofpacket                                                                       : std_logic;                      -- id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal id_router_001_src_data                                                                                : std_logic_vector(99 downto 0);  -- id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	signal id_router_001_src_channel                                                                             : std_logic_vector(3 downto 0);   -- id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	signal id_router_001_src_ready                                                                               : std_logic;                      -- rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	signal cmd_xbar_demux_src2_ready                                                                             : std_logic;                      -- cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src2_ready
	signal id_router_002_src_endofpacket                                                                         : std_logic;                      -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                               : std_logic;                      -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                                       : std_logic;                      -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                                : std_logic_vector(99 downto 0);  -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                             : std_logic_vector(3 downto 0);   -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                               : std_logic;                      -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal cmd_xbar_mux_003_src_endofpacket                                                                      : std_logic;                      -- cmd_xbar_mux_003:src_endofpacket -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_003_src_valid                                                                            : std_logic;                      -- cmd_xbar_mux_003:src_valid -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_003_src_startofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_003:src_startofpacket -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_003_src_data                                                                             : std_logic_vector(99 downto 0);  -- cmd_xbar_mux_003:src_data -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_003_src_channel                                                                          : std_logic_vector(3 downto 0);   -- cmd_xbar_mux_003:src_channel -> cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_003_src_ready                                                                            : std_logic;                      -- cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	signal id_router_003_src_endofpacket                                                                         : std_logic;                      -- id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal id_router_003_src_valid                                                                               : std_logic;                      -- id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	signal id_router_003_src_startofpacket                                                                       : std_logic;                      -- id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal id_router_003_src_data                                                                                : std_logic_vector(99 downto 0);  -- id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	signal id_router_003_src_channel                                                                             : std_logic_vector(3 downto 0);   -- id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	signal id_router_003_src_ready                                                                               : std_logic;                      -- rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	signal cmd_xbar_demux_002_src0_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	signal cmd_xbar_demux_002_src0_valid                                                                         : std_logic;                      -- cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_004:sink0_valid
	signal cmd_xbar_demux_002_src0_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	signal cmd_xbar_demux_002_src0_data                                                                          : std_logic_vector(100 downto 0); -- cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_004:sink0_data
	signal cmd_xbar_demux_002_src0_channel                                                                       : std_logic_vector(3 downto 0);   -- cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_004:sink0_channel
	signal cmd_xbar_demux_002_src0_ready                                                                         : std_logic;                      -- cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux_002:src0_ready
	signal cmd_xbar_demux_003_src0_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	signal cmd_xbar_demux_003_src0_valid                                                                         : std_logic;                      -- cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_004:sink1_valid
	signal cmd_xbar_demux_003_src0_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	signal cmd_xbar_demux_003_src0_data                                                                          : std_logic_vector(100 downto 0); -- cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_004:sink1_data
	signal cmd_xbar_demux_003_src0_channel                                                                       : std_logic_vector(3 downto 0);   -- cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_004:sink1_channel
	signal cmd_xbar_demux_003_src0_ready                                                                         : std_logic;                      -- cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_003:src0_ready
	signal cmd_xbar_demux_004_src0_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_004:sink2_endofpacket
	signal cmd_xbar_demux_004_src0_valid                                                                         : std_logic;                      -- cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_004:sink2_valid
	signal cmd_xbar_demux_004_src0_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_004:sink2_startofpacket
	signal cmd_xbar_demux_004_src0_data                                                                          : std_logic_vector(100 downto 0); -- cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_004:sink2_data
	signal cmd_xbar_demux_004_src0_channel                                                                       : std_logic_vector(3 downto 0);   -- cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_004:sink2_channel
	signal cmd_xbar_demux_004_src0_ready                                                                         : std_logic;                      -- cmd_xbar_mux_004:sink2_ready -> cmd_xbar_demux_004:src0_ready
	signal cmd_xbar_demux_005_src0_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_005:src0_endofpacket -> cmd_xbar_mux_004:sink3_endofpacket
	signal cmd_xbar_demux_005_src0_valid                                                                         : std_logic;                      -- cmd_xbar_demux_005:src0_valid -> cmd_xbar_mux_004:sink3_valid
	signal cmd_xbar_demux_005_src0_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_005:src0_startofpacket -> cmd_xbar_mux_004:sink3_startofpacket
	signal cmd_xbar_demux_005_src0_data                                                                          : std_logic_vector(100 downto 0); -- cmd_xbar_demux_005:src0_data -> cmd_xbar_mux_004:sink3_data
	signal cmd_xbar_demux_005_src0_channel                                                                       : std_logic_vector(3 downto 0);   -- cmd_xbar_demux_005:src0_channel -> cmd_xbar_mux_004:sink3_channel
	signal cmd_xbar_demux_005_src0_ready                                                                         : std_logic;                      -- cmd_xbar_mux_004:sink3_ready -> cmd_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_004:src0_endofpacket -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_004:src0_valid -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_004:src0_startofpacket -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                          : std_logic_vector(100 downto 0); -- rsp_xbar_demux_004:src0_data -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_demux_004_src0_channel                                                                       : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_004:src0_channel -> sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_demux_004_src1_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_004:src1_endofpacket -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_demux_004_src1_valid                                                                         : std_logic;                      -- rsp_xbar_demux_004:src1_valid -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_demux_004_src1_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_004:src1_startofpacket -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_demux_004_src1_data                                                                          : std_logic_vector(100 downto 0); -- rsp_xbar_demux_004:src1_data -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_demux_004_src1_channel                                                                       : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_004:src1_channel -> sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_demux_004_src2_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_004:src2_endofpacket -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_demux_004_src2_valid                                                                         : std_logic;                      -- rsp_xbar_demux_004:src2_valid -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_demux_004_src2_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_004:src2_startofpacket -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_demux_004_src2_data                                                                          : std_logic_vector(100 downto 0); -- rsp_xbar_demux_004:src2_data -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_demux_004_src2_channel                                                                       : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_004:src2_channel -> sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_demux_004_src3_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_004:src3_endofpacket -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_demux_004_src3_valid                                                                         : std_logic;                      -- rsp_xbar_demux_004:src3_valid -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_demux_004_src3_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_004:src3_startofpacket -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_demux_004_src3_data                                                                          : std_logic_vector(100 downto 0); -- rsp_xbar_demux_004:src3_data -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_demux_004_src3_channel                                                                       : std_logic_vector(3 downto 0);   -- rsp_xbar_demux_004:src3_channel -> sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_channel
	signal addr_router_002_src_endofpacket                                                                       : std_logic;                      -- addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	signal addr_router_002_src_valid                                                                             : std_logic;                      -- addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	signal addr_router_002_src_startofpacket                                                                     : std_logic;                      -- addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	signal addr_router_002_src_data                                                                              : std_logic_vector(100 downto 0); -- addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	signal addr_router_002_src_channel                                                                           : std_logic_vector(3 downto 0);   -- addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	signal addr_router_002_src_ready                                                                             : std_logic;                      -- cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	signal rsp_xbar_demux_004_src0_ready                                                                         : std_logic;                      -- sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_004:src0_ready
	signal addr_router_003_src_endofpacket                                                                       : std_logic;                      -- addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	signal addr_router_003_src_valid                                                                             : std_logic;                      -- addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	signal addr_router_003_src_startofpacket                                                                     : std_logic;                      -- addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	signal addr_router_003_src_data                                                                              : std_logic_vector(100 downto 0); -- addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	signal addr_router_003_src_channel                                                                           : std_logic_vector(3 downto 0);   -- addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	signal addr_router_003_src_ready                                                                             : std_logic;                      -- cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	signal rsp_xbar_demux_004_src1_ready                                                                         : std_logic;                      -- sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_004:src1_ready
	signal addr_router_004_src_endofpacket                                                                       : std_logic;                      -- addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	signal addr_router_004_src_valid                                                                             : std_logic;                      -- addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	signal addr_router_004_src_startofpacket                                                                     : std_logic;                      -- addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	signal addr_router_004_src_data                                                                              : std_logic_vector(100 downto 0); -- addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	signal addr_router_004_src_channel                                                                           : std_logic_vector(3 downto 0);   -- addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	signal addr_router_004_src_ready                                                                             : std_logic;                      -- cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	signal rsp_xbar_demux_004_src2_ready                                                                         : std_logic;                      -- sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_004:src2_ready
	signal addr_router_005_src_endofpacket                                                                       : std_logic;                      -- addr_router_005:src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	signal addr_router_005_src_valid                                                                             : std_logic;                      -- addr_router_005:src_valid -> cmd_xbar_demux_005:sink_valid
	signal addr_router_005_src_startofpacket                                                                     : std_logic;                      -- addr_router_005:src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	signal addr_router_005_src_data                                                                              : std_logic_vector(100 downto 0); -- addr_router_005:src_data -> cmd_xbar_demux_005:sink_data
	signal addr_router_005_src_channel                                                                           : std_logic_vector(3 downto 0);   -- addr_router_005:src_channel -> cmd_xbar_demux_005:sink_channel
	signal addr_router_005_src_ready                                                                             : std_logic;                      -- cmd_xbar_demux_005:sink_ready -> addr_router_005:src_ready
	signal rsp_xbar_demux_004_src3_ready                                                                         : std_logic;                      -- sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_004:src3_ready
	signal cmd_xbar_mux_004_src_endofpacket                                                                      : std_logic;                      -- cmd_xbar_mux_004:src_endofpacket -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_004_src_valid                                                                            : std_logic;                      -- cmd_xbar_mux_004:src_valid -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_004_src_startofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_004:src_startofpacket -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_004_src_data                                                                             : std_logic_vector(100 downto 0); -- cmd_xbar_mux_004:src_data -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_004_src_channel                                                                          : std_logic_vector(3 downto 0);   -- cmd_xbar_mux_004:src_channel -> dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_004_src_ready                                                                            : std_logic;                      -- dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	signal id_router_004_src_endofpacket                                                                         : std_logic;                      -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                               : std_logic;                      -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                       : std_logic;                      -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                                : std_logic_vector(100 downto 0); -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                             : std_logic_vector(3 downto 0);   -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                               : std_logic;                      -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_demux_006_src0_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_006:src0_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	signal cmd_xbar_demux_006_src0_valid                                                                         : std_logic;                      -- cmd_xbar_demux_006:src0_valid -> cmd_xbar_mux_005:sink0_valid
	signal cmd_xbar_demux_006_src0_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_006:src0_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	signal cmd_xbar_demux_006_src0_data                                                                          : std_logic_vector(93 downto 0);  -- cmd_xbar_demux_006:src0_data -> cmd_xbar_mux_005:sink0_data
	signal cmd_xbar_demux_006_src0_channel                                                                       : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_006:src0_channel -> cmd_xbar_mux_005:sink0_channel
	signal cmd_xbar_demux_006_src0_ready                                                                         : std_logic;                      -- cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux_006:src0_ready
	signal cmd_xbar_demux_007_src0_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_007:src0_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	signal cmd_xbar_demux_007_src0_valid                                                                         : std_logic;                      -- cmd_xbar_demux_007:src0_valid -> cmd_xbar_mux_005:sink1_valid
	signal cmd_xbar_demux_007_src0_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_007:src0_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	signal cmd_xbar_demux_007_src0_data                                                                          : std_logic_vector(93 downto 0);  -- cmd_xbar_demux_007:src0_data -> cmd_xbar_mux_005:sink1_data
	signal cmd_xbar_demux_007_src0_channel                                                                       : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_007:src0_channel -> cmd_xbar_mux_005:sink1_channel
	signal cmd_xbar_demux_007_src0_ready                                                                         : std_logic;                      -- cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_007:src0_ready
	signal cmd_xbar_demux_007_src1_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_007:src1_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_007_src1_valid                                                                         : std_logic;                      -- cmd_xbar_demux_007:src1_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_007_src1_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_007:src1_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_007_src1_data                                                                          : std_logic_vector(93 downto 0);  -- cmd_xbar_demux_007:src1_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_007_src1_channel                                                                       : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_007:src1_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_007_src2_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_007:src2_endofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_007_src2_valid                                                                         : std_logic;                      -- cmd_xbar_demux_007:src2_valid -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_007_src2_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_007:src2_startofpacket -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_007_src2_data                                                                          : std_logic_vector(93 downto 0);  -- cmd_xbar_demux_007:src2_data -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_007_src2_channel                                                                       : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_007:src2_channel -> tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_007_src3_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_007:src3_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_007_src3_valid                                                                         : std_logic;                      -- cmd_xbar_demux_007:src3_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_007_src3_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_007:src3_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_007_src3_data                                                                          : std_logic_vector(93 downto 0);  -- cmd_xbar_demux_007:src3_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_007_src3_channel                                                                       : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_007:src3_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_007_src4_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_007:src4_endofpacket -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_007_src4_valid                                                                         : std_logic;                      -- cmd_xbar_demux_007:src4_valid -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_007_src4_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_007:src4_startofpacket -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_007_src4_data                                                                          : std_logic_vector(93 downto 0);  -- cmd_xbar_demux_007:src4_data -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_007_src4_channel                                                                       : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_007:src4_channel -> linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_007_src5_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_007:src5_endofpacket -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_007_src5_valid                                                                         : std_logic;                      -- cmd_xbar_demux_007:src5_valid -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_007_src5_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_007:src5_startofpacket -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_007_src5_data                                                                          : std_logic_vector(93 downto 0);  -- cmd_xbar_demux_007:src5_data -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_007_src5_channel                                                                       : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_007:src5_channel -> gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_007_src6_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_007:src6_endofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_007_src6_valid                                                                         : std_logic;                      -- cmd_xbar_demux_007:src6_valid -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_007_src6_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_007:src6_startofpacket -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_007_src6_data                                                                          : std_logic_vector(93 downto 0);  -- cmd_xbar_demux_007:src6_data -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_007_src6_channel                                                                       : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_007:src6_channel -> sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_007_src7_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_007:src7_endofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_007_src7_valid                                                                         : std_logic;                      -- cmd_xbar_demux_007:src7_valid -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_007_src7_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_007:src7_startofpacket -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_007_src7_data                                                                          : std_logic_vector(93 downto 0);  -- cmd_xbar_demux_007:src7_data -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_007_src7_channel                                                                       : std_logic_vector(7 downto 0);   -- cmd_xbar_demux_007:src7_channel -> sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_channel
	signal rsp_xbar_demux_005_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_005:src0_endofpacket -> dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_005:src0_valid -> dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_005:src0_startofpacket -> dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                          : std_logic_vector(93 downto 0);  -- rsp_xbar_demux_005:src0_data -> dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_demux_005_src0_channel                                                                       : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_005:src0_channel -> dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_demux_005_src1_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_007:sink0_endofpacket
	signal rsp_xbar_demux_005_src1_valid                                                                         : std_logic;                      -- rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_007:sink0_valid
	signal rsp_xbar_demux_005_src1_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_007:sink0_startofpacket
	signal rsp_xbar_demux_005_src1_data                                                                          : std_logic_vector(93 downto 0);  -- rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_007:sink0_data
	signal rsp_xbar_demux_005_src1_channel                                                                       : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_007:sink0_channel
	signal rsp_xbar_demux_005_src1_ready                                                                         : std_logic;                      -- rsp_xbar_mux_007:sink0_ready -> rsp_xbar_demux_005:src1_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_007:sink1_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_007:sink1_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_007:sink1_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                          : std_logic_vector(93 downto 0);  -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_007:sink1_data
	signal rsp_xbar_demux_006_src0_channel                                                                       : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_007:sink1_channel
	signal rsp_xbar_demux_006_src0_ready                                                                         : std_logic;                      -- rsp_xbar_mux_007:sink1_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_007:sink2_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_007:sink2_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_007:sink2_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                          : std_logic_vector(93 downto 0);  -- rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_007:sink2_data
	signal rsp_xbar_demux_007_src0_channel                                                                       : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_007:sink2_channel
	signal rsp_xbar_demux_007_src0_ready                                                                         : std_logic;                      -- rsp_xbar_mux_007:sink2_ready -> rsp_xbar_demux_007:src0_ready
	signal rsp_xbar_demux_008_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_007:sink3_endofpacket
	signal rsp_xbar_demux_008_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_007:sink3_valid
	signal rsp_xbar_demux_008_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_007:sink3_startofpacket
	signal rsp_xbar_demux_008_src0_data                                                                          : std_logic_vector(93 downto 0);  -- rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_007:sink3_data
	signal rsp_xbar_demux_008_src0_channel                                                                       : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_007:sink3_channel
	signal rsp_xbar_demux_008_src0_ready                                                                         : std_logic;                      -- rsp_xbar_mux_007:sink3_ready -> rsp_xbar_demux_008:src0_ready
	signal rsp_xbar_demux_009_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_007:sink4_endofpacket
	signal rsp_xbar_demux_009_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_007:sink4_valid
	signal rsp_xbar_demux_009_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_007:sink4_startofpacket
	signal rsp_xbar_demux_009_src0_data                                                                          : std_logic_vector(93 downto 0);  -- rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_007:sink4_data
	signal rsp_xbar_demux_009_src0_channel                                                                       : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_007:sink4_channel
	signal rsp_xbar_demux_009_src0_ready                                                                         : std_logic;                      -- rsp_xbar_mux_007:sink4_ready -> rsp_xbar_demux_009:src0_ready
	signal rsp_xbar_demux_010_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_007:sink5_endofpacket
	signal rsp_xbar_demux_010_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_007:sink5_valid
	signal rsp_xbar_demux_010_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_007:sink5_startofpacket
	signal rsp_xbar_demux_010_src0_data                                                                          : std_logic_vector(93 downto 0);  -- rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_007:sink5_data
	signal rsp_xbar_demux_010_src0_channel                                                                       : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_007:sink5_channel
	signal rsp_xbar_demux_010_src0_ready                                                                         : std_logic;                      -- rsp_xbar_mux_007:sink5_ready -> rsp_xbar_demux_010:src0_ready
	signal rsp_xbar_demux_011_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_007:sink6_endofpacket
	signal rsp_xbar_demux_011_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_007:sink6_valid
	signal rsp_xbar_demux_011_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_007:sink6_startofpacket
	signal rsp_xbar_demux_011_src0_data                                                                          : std_logic_vector(93 downto 0);  -- rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_007:sink6_data
	signal rsp_xbar_demux_011_src0_channel                                                                       : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_007:sink6_channel
	signal rsp_xbar_demux_011_src0_ready                                                                         : std_logic;                      -- rsp_xbar_mux_007:sink6_ready -> rsp_xbar_demux_011:src0_ready
	signal rsp_xbar_demux_012_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_007:sink7_endofpacket
	signal rsp_xbar_demux_012_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_007:sink7_valid
	signal rsp_xbar_demux_012_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_007:sink7_startofpacket
	signal rsp_xbar_demux_012_src0_data                                                                          : std_logic_vector(93 downto 0);  -- rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_007:sink7_data
	signal rsp_xbar_demux_012_src0_channel                                                                       : std_logic_vector(7 downto 0);   -- rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_007:sink7_channel
	signal rsp_xbar_demux_012_src0_ready                                                                         : std_logic;                      -- rsp_xbar_mux_007:sink7_ready -> rsp_xbar_demux_012:src0_ready
	signal addr_router_006_src_endofpacket                                                                       : std_logic;                      -- addr_router_006:src_endofpacket -> cmd_xbar_demux_006:sink_endofpacket
	signal addr_router_006_src_valid                                                                             : std_logic;                      -- addr_router_006:src_valid -> cmd_xbar_demux_006:sink_valid
	signal addr_router_006_src_startofpacket                                                                     : std_logic;                      -- addr_router_006:src_startofpacket -> cmd_xbar_demux_006:sink_startofpacket
	signal addr_router_006_src_data                                                                              : std_logic_vector(93 downto 0);  -- addr_router_006:src_data -> cmd_xbar_demux_006:sink_data
	signal addr_router_006_src_channel                                                                           : std_logic_vector(7 downto 0);   -- addr_router_006:src_channel -> cmd_xbar_demux_006:sink_channel
	signal addr_router_006_src_ready                                                                             : std_logic;                      -- cmd_xbar_demux_006:sink_ready -> addr_router_006:src_ready
	signal rsp_xbar_demux_005_src0_ready                                                                         : std_logic;                      -- dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_005:src0_ready
	signal limiter_002_cmd_src_endofpacket                                                                       : std_logic;                      -- limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_007:sink_endofpacket
	signal limiter_002_cmd_src_startofpacket                                                                     : std_logic;                      -- limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_007:sink_startofpacket
	signal limiter_002_cmd_src_data                                                                              : std_logic_vector(93 downto 0);  -- limiter_002:cmd_src_data -> cmd_xbar_demux_007:sink_data
	signal limiter_002_cmd_src_channel                                                                           : std_logic_vector(7 downto 0);   -- limiter_002:cmd_src_channel -> cmd_xbar_demux_007:sink_channel
	signal limiter_002_cmd_src_ready                                                                             : std_logic;                      -- cmd_xbar_demux_007:sink_ready -> limiter_002:cmd_src_ready
	signal rsp_xbar_mux_007_src_endofpacket                                                                      : std_logic;                      -- rsp_xbar_mux_007:src_endofpacket -> limiter_002:rsp_sink_endofpacket
	signal rsp_xbar_mux_007_src_valid                                                                            : std_logic;                      -- rsp_xbar_mux_007:src_valid -> limiter_002:rsp_sink_valid
	signal rsp_xbar_mux_007_src_startofpacket                                                                    : std_logic;                      -- rsp_xbar_mux_007:src_startofpacket -> limiter_002:rsp_sink_startofpacket
	signal rsp_xbar_mux_007_src_data                                                                             : std_logic_vector(93 downto 0);  -- rsp_xbar_mux_007:src_data -> limiter_002:rsp_sink_data
	signal rsp_xbar_mux_007_src_channel                                                                          : std_logic_vector(7 downto 0);   -- rsp_xbar_mux_007:src_channel -> limiter_002:rsp_sink_channel
	signal rsp_xbar_mux_007_src_ready                                                                            : std_logic;                      -- limiter_002:rsp_sink_ready -> rsp_xbar_mux_007:src_ready
	signal cmd_xbar_mux_005_src_endofpacket                                                                      : std_logic;                      -- cmd_xbar_mux_005:src_endofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_005_src_valid                                                                            : std_logic;                      -- cmd_xbar_mux_005:src_valid -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_005_src_startofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_005:src_startofpacket -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_005_src_data                                                                             : std_logic_vector(93 downto 0);  -- cmd_xbar_mux_005:src_data -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_005_src_channel                                                                          : std_logic_vector(7 downto 0);   -- cmd_xbar_mux_005:src_channel -> descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_005_src_ready                                                                            : std_logic;                      -- descriptor_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	signal id_router_005_src_endofpacket                                                                         : std_logic;                      -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                               : std_logic;                      -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                       : std_logic;                      -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                                : std_logic_vector(93 downto 0);  -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                             : std_logic_vector(7 downto 0);   -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                               : std_logic;                      -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_demux_007_src1_ready                                                                         : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src1_ready
	signal id_router_006_src_endofpacket                                                                         : std_logic;                      -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                               : std_logic;                      -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                       : std_logic;                      -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                                : std_logic_vector(93 downto 0);  -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                             : std_logic_vector(7 downto 0);   -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                               : std_logic;                      -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_demux_007_src2_ready                                                                         : std_logic;                      -- tse_mac_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src2_ready
	signal id_router_007_src_endofpacket                                                                         : std_logic;                      -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                               : std_logic;                      -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                                       : std_logic;                      -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                                : std_logic_vector(93 downto 0);  -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                             : std_logic_vector(7 downto 0);   -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                               : std_logic;                      -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal cmd_xbar_demux_007_src3_ready                                                                         : std_logic;                      -- sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src3_ready
	signal id_router_008_src_endofpacket                                                                         : std_logic;                      -- id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	signal id_router_008_src_valid                                                                               : std_logic;                      -- id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	signal id_router_008_src_startofpacket                                                                       : std_logic;                      -- id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	signal id_router_008_src_data                                                                                : std_logic_vector(93 downto 0);  -- id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	signal id_router_008_src_channel                                                                             : std_logic_vector(7 downto 0);   -- id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	signal id_router_008_src_ready                                                                               : std_logic;                      -- rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	signal cmd_xbar_demux_007_src4_ready                                                                         : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src4_ready
	signal id_router_009_src_endofpacket                                                                         : std_logic;                      -- id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	signal id_router_009_src_valid                                                                               : std_logic;                      -- id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	signal id_router_009_src_startofpacket                                                                       : std_logic;                      -- id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	signal id_router_009_src_data                                                                                : std_logic_vector(93 downto 0);  -- id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	signal id_router_009_src_channel                                                                             : std_logic_vector(7 downto 0);   -- id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	signal id_router_009_src_ready                                                                               : std_logic;                      -- rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	signal cmd_xbar_demux_007_src5_ready                                                                         : std_logic;                      -- gtp_regif_0_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src5_ready
	signal id_router_010_src_endofpacket                                                                         : std_logic;                      -- id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	signal id_router_010_src_valid                                                                               : std_logic;                      -- id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	signal id_router_010_src_startofpacket                                                                       : std_logic;                      -- id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	signal id_router_010_src_data                                                                                : std_logic_vector(93 downto 0);  -- id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	signal id_router_010_src_channel                                                                             : std_logic_vector(7 downto 0);   -- id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	signal id_router_010_src_ready                                                                               : std_logic;                      -- rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	signal cmd_xbar_demux_007_src6_ready                                                                         : std_logic;                      -- sgdma_tx_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src6_ready
	signal id_router_011_src_endofpacket                                                                         : std_logic;                      -- id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	signal id_router_011_src_valid                                                                               : std_logic;                      -- id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	signal id_router_011_src_startofpacket                                                                       : std_logic;                      -- id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	signal id_router_011_src_data                                                                                : std_logic_vector(93 downto 0);  -- id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	signal id_router_011_src_channel                                                                             : std_logic_vector(7 downto 0);   -- id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	signal id_router_011_src_ready                                                                               : std_logic;                      -- rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	signal cmd_xbar_demux_007_src7_ready                                                                         : std_logic;                      -- sgdma_rx_csr_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src7_ready
	signal id_router_012_src_endofpacket                                                                         : std_logic;                      -- id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	signal id_router_012_src_valid                                                                               : std_logic;                      -- id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	signal id_router_012_src_startofpacket                                                                       : std_logic;                      -- id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	signal id_router_012_src_data                                                                                : std_logic_vector(93 downto 0);  -- id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	signal id_router_012_src_channel                                                                             : std_logic_vector(7 downto 0);   -- id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	signal id_router_012_src_ready                                                                               : std_logic;                      -- rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	signal cmd_xbar_demux_008_src0_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_008:src0_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_demux_008_src0_valid                                                                         : std_logic;                      -- cmd_xbar_demux_008:src0_valid -> width_adapter:in_valid
	signal cmd_xbar_demux_008_src0_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_008:src0_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_demux_008_src0_data                                                                          : std_logic_vector(94 downto 0);  -- cmd_xbar_demux_008:src0_data -> width_adapter:in_data
	signal cmd_xbar_demux_008_src0_channel                                                                       : std_logic_vector(1 downto 0);   -- cmd_xbar_demux_008:src0_channel -> width_adapter:in_channel
	signal cmd_xbar_demux_008_src1_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_008:src1_endofpacket -> width_adapter_002:in_endofpacket
	signal cmd_xbar_demux_008_src1_valid                                                                         : std_logic;                      -- cmd_xbar_demux_008:src1_valid -> width_adapter_002:in_valid
	signal cmd_xbar_demux_008_src1_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_008:src1_startofpacket -> width_adapter_002:in_startofpacket
	signal cmd_xbar_demux_008_src1_data                                                                          : std_logic_vector(94 downto 0);  -- cmd_xbar_demux_008:src1_data -> width_adapter_002:in_data
	signal cmd_xbar_demux_008_src1_channel                                                                       : std_logic_vector(1 downto 0);   -- cmd_xbar_demux_008:src1_channel -> width_adapter_002:in_channel
	signal rsp_xbar_demux_013_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_008:sink0_endofpacket
	signal rsp_xbar_demux_013_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_008:sink0_valid
	signal rsp_xbar_demux_013_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_008:sink0_startofpacket
	signal rsp_xbar_demux_013_src0_data                                                                          : std_logic_vector(94 downto 0);  -- rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_008:sink0_data
	signal rsp_xbar_demux_013_src0_channel                                                                       : std_logic_vector(1 downto 0);   -- rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_008:sink0_channel
	signal rsp_xbar_demux_013_src0_ready                                                                         : std_logic;                      -- rsp_xbar_mux_008:sink0_ready -> rsp_xbar_demux_013:src0_ready
	signal rsp_xbar_demux_014_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_008:sink1_endofpacket
	signal rsp_xbar_demux_014_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_008:sink1_valid
	signal rsp_xbar_demux_014_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_008:sink1_startofpacket
	signal rsp_xbar_demux_014_src0_data                                                                          : std_logic_vector(94 downto 0);  -- rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_008:sink1_data
	signal rsp_xbar_demux_014_src0_channel                                                                       : std_logic_vector(1 downto 0);   -- rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_008:sink1_channel
	signal rsp_xbar_demux_014_src0_ready                                                                         : std_logic;                      -- rsp_xbar_mux_008:sink1_ready -> rsp_xbar_demux_014:src0_ready
	signal limiter_003_cmd_src_endofpacket                                                                       : std_logic;                      -- limiter_003:cmd_src_endofpacket -> cmd_xbar_demux_008:sink_endofpacket
	signal limiter_003_cmd_src_startofpacket                                                                     : std_logic;                      -- limiter_003:cmd_src_startofpacket -> cmd_xbar_demux_008:sink_startofpacket
	signal limiter_003_cmd_src_data                                                                              : std_logic_vector(94 downto 0);  -- limiter_003:cmd_src_data -> cmd_xbar_demux_008:sink_data
	signal limiter_003_cmd_src_channel                                                                           : std_logic_vector(1 downto 0);   -- limiter_003:cmd_src_channel -> cmd_xbar_demux_008:sink_channel
	signal limiter_003_cmd_src_ready                                                                             : std_logic;                      -- cmd_xbar_demux_008:sink_ready -> limiter_003:cmd_src_ready
	signal rsp_xbar_mux_008_src_endofpacket                                                                      : std_logic;                      -- rsp_xbar_mux_008:src_endofpacket -> limiter_003:rsp_sink_endofpacket
	signal rsp_xbar_mux_008_src_valid                                                                            : std_logic;                      -- rsp_xbar_mux_008:src_valid -> limiter_003:rsp_sink_valid
	signal rsp_xbar_mux_008_src_startofpacket                                                                    : std_logic;                      -- rsp_xbar_mux_008:src_startofpacket -> limiter_003:rsp_sink_startofpacket
	signal rsp_xbar_mux_008_src_data                                                                             : std_logic_vector(94 downto 0);  -- rsp_xbar_mux_008:src_data -> limiter_003:rsp_sink_data
	signal rsp_xbar_mux_008_src_channel                                                                          : std_logic_vector(1 downto 0);   -- rsp_xbar_mux_008:src_channel -> limiter_003:rsp_sink_channel
	signal rsp_xbar_mux_008_src_ready                                                                            : std_logic;                      -- limiter_003:rsp_sink_ready -> rsp_xbar_mux_008:src_ready
	signal cmd_xbar_demux_009_src0_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_009:src0_endofpacket -> cmd_xbar_mux_015:sink0_endofpacket
	signal cmd_xbar_demux_009_src0_valid                                                                         : std_logic;                      -- cmd_xbar_demux_009:src0_valid -> cmd_xbar_mux_015:sink0_valid
	signal cmd_xbar_demux_009_src0_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_009:src0_startofpacket -> cmd_xbar_mux_015:sink0_startofpacket
	signal cmd_xbar_demux_009_src0_data                                                                          : std_logic_vector(98 downto 0);  -- cmd_xbar_demux_009:src0_data -> cmd_xbar_mux_015:sink0_data
	signal cmd_xbar_demux_009_src0_channel                                                                       : std_logic_vector(1 downto 0);   -- cmd_xbar_demux_009:src0_channel -> cmd_xbar_mux_015:sink0_channel
	signal cmd_xbar_demux_009_src0_ready                                                                         : std_logic;                      -- cmd_xbar_mux_015:sink0_ready -> cmd_xbar_demux_009:src0_ready
	signal cmd_xbar_demux_010_src0_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_010:src0_endofpacket -> cmd_xbar_mux_015:sink1_endofpacket
	signal cmd_xbar_demux_010_src0_valid                                                                         : std_logic;                      -- cmd_xbar_demux_010:src0_valid -> cmd_xbar_mux_015:sink1_valid
	signal cmd_xbar_demux_010_src0_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_010:src0_startofpacket -> cmd_xbar_mux_015:sink1_startofpacket
	signal cmd_xbar_demux_010_src0_data                                                                          : std_logic_vector(98 downto 0);  -- cmd_xbar_demux_010:src0_data -> cmd_xbar_mux_015:sink1_data
	signal cmd_xbar_demux_010_src0_channel                                                                       : std_logic_vector(1 downto 0);   -- cmd_xbar_demux_010:src0_channel -> cmd_xbar_mux_015:sink1_channel
	signal cmd_xbar_demux_010_src0_ready                                                                         : std_logic;                      -- cmd_xbar_mux_015:sink1_ready -> cmd_xbar_demux_010:src0_ready
	signal rsp_xbar_demux_015_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_015:src0_endofpacket -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_demux_015_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_015:src0_valid -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_demux_015_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_015:src0_startofpacket -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_demux_015_src0_data                                                                          : std_logic_vector(98 downto 0);  -- rsp_xbar_demux_015:src0_data -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_demux_015_src0_channel                                                                       : std_logic_vector(1 downto 0);   -- rsp_xbar_demux_015:src0_channel -> sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_demux_015_src1_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_015:src1_endofpacket -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_demux_015_src1_valid                                                                         : std_logic;                      -- rsp_xbar_demux_015:src1_valid -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_demux_015_src1_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_015:src1_startofpacket -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_demux_015_src1_data                                                                          : std_logic_vector(98 downto 0);  -- rsp_xbar_demux_015:src1_data -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_demux_015_src1_channel                                                                       : std_logic_vector(1 downto 0);   -- rsp_xbar_demux_015:src1_channel -> sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_channel
	signal addr_router_009_src_endofpacket                                                                       : std_logic;                      -- addr_router_009:src_endofpacket -> cmd_xbar_demux_009:sink_endofpacket
	signal addr_router_009_src_valid                                                                             : std_logic;                      -- addr_router_009:src_valid -> cmd_xbar_demux_009:sink_valid
	signal addr_router_009_src_startofpacket                                                                     : std_logic;                      -- addr_router_009:src_startofpacket -> cmd_xbar_demux_009:sink_startofpacket
	signal addr_router_009_src_data                                                                              : std_logic_vector(98 downto 0);  -- addr_router_009:src_data -> cmd_xbar_demux_009:sink_data
	signal addr_router_009_src_channel                                                                           : std_logic_vector(1 downto 0);   -- addr_router_009:src_channel -> cmd_xbar_demux_009:sink_channel
	signal addr_router_009_src_ready                                                                             : std_logic;                      -- cmd_xbar_demux_009:sink_ready -> addr_router_009:src_ready
	signal rsp_xbar_demux_015_src0_ready                                                                         : std_logic;                      -- sgdma_tx_m_read_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_015:src0_ready
	signal addr_router_010_src_endofpacket                                                                       : std_logic;                      -- addr_router_010:src_endofpacket -> cmd_xbar_demux_010:sink_endofpacket
	signal addr_router_010_src_valid                                                                             : std_logic;                      -- addr_router_010:src_valid -> cmd_xbar_demux_010:sink_valid
	signal addr_router_010_src_startofpacket                                                                     : std_logic;                      -- addr_router_010:src_startofpacket -> cmd_xbar_demux_010:sink_startofpacket
	signal addr_router_010_src_data                                                                              : std_logic_vector(98 downto 0);  -- addr_router_010:src_data -> cmd_xbar_demux_010:sink_data
	signal addr_router_010_src_channel                                                                           : std_logic_vector(1 downto 0);   -- addr_router_010:src_channel -> cmd_xbar_demux_010:sink_channel
	signal addr_router_010_src_ready                                                                             : std_logic;                      -- cmd_xbar_demux_010:sink_ready -> addr_router_010:src_ready
	signal rsp_xbar_demux_015_src1_ready                                                                         : std_logic;                      -- sgdma_rx_m_write_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_015:src1_ready
	signal cmd_xbar_mux_015_src_endofpacket                                                                      : std_logic;                      -- cmd_xbar_mux_015:src_endofpacket -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_015_src_valid                                                                            : std_logic;                      -- cmd_xbar_mux_015:src_valid -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_015_src_startofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_015:src_startofpacket -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_015_src_data                                                                             : std_logic_vector(98 downto 0);  -- cmd_xbar_mux_015:src_data -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_015_src_channel                                                                          : std_logic_vector(1 downto 0);   -- cmd_xbar_mux_015:src_channel -> tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_015_src_ready                                                                            : std_logic;                      -- tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_015:src_ready
	signal id_router_015_src_endofpacket                                                                         : std_logic;                      -- id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	signal id_router_015_src_valid                                                                               : std_logic;                      -- id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	signal id_router_015_src_startofpacket                                                                       : std_logic;                      -- id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	signal id_router_015_src_data                                                                                : std_logic_vector(98 downto 0);  -- id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	signal id_router_015_src_channel                                                                             : std_logic_vector(1 downto 0);   -- id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	signal id_router_015_src_ready                                                                               : std_logic;                      -- rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	signal cmd_xbar_demux_011_src0_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_011:src0_endofpacket -> cmd_xbar_mux_016:sink0_endofpacket
	signal cmd_xbar_demux_011_src0_valid                                                                         : std_logic;                      -- cmd_xbar_demux_011:src0_valid -> cmd_xbar_mux_016:sink0_valid
	signal cmd_xbar_demux_011_src0_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_011:src0_startofpacket -> cmd_xbar_mux_016:sink0_startofpacket
	signal cmd_xbar_demux_011_src0_data                                                                          : std_logic_vector(96 downto 0);  -- cmd_xbar_demux_011:src0_data -> cmd_xbar_mux_016:sink0_data
	signal cmd_xbar_demux_011_src0_channel                                                                       : std_logic_vector(1 downto 0);   -- cmd_xbar_demux_011:src0_channel -> cmd_xbar_mux_016:sink0_channel
	signal cmd_xbar_demux_011_src0_ready                                                                         : std_logic;                      -- cmd_xbar_mux_016:sink0_ready -> cmd_xbar_demux_011:src0_ready
	signal cmd_xbar_demux_012_src0_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_012:src0_endofpacket -> cmd_xbar_mux_016:sink1_endofpacket
	signal cmd_xbar_demux_012_src0_valid                                                                         : std_logic;                      -- cmd_xbar_demux_012:src0_valid -> cmd_xbar_mux_016:sink1_valid
	signal cmd_xbar_demux_012_src0_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_012:src0_startofpacket -> cmd_xbar_mux_016:sink1_startofpacket
	signal cmd_xbar_demux_012_src0_data                                                                          : std_logic_vector(96 downto 0);  -- cmd_xbar_demux_012:src0_data -> cmd_xbar_mux_016:sink1_data
	signal cmd_xbar_demux_012_src0_channel                                                                       : std_logic_vector(1 downto 0);   -- cmd_xbar_demux_012:src0_channel -> cmd_xbar_mux_016:sink1_channel
	signal cmd_xbar_demux_012_src0_ready                                                                         : std_logic;                      -- cmd_xbar_mux_016:sink1_ready -> cmd_xbar_demux_012:src0_ready
	signal rsp_xbar_demux_016_src0_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_016:src0_endofpacket -> tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_demux_016_src0_valid                                                                         : std_logic;                      -- rsp_xbar_demux_016:src0_valid -> tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_demux_016_src0_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_016:src0_startofpacket -> tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_demux_016_src0_data                                                                          : std_logic_vector(96 downto 0);  -- rsp_xbar_demux_016:src0_data -> tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_demux_016_src0_channel                                                                       : std_logic_vector(1 downto 0);   -- rsp_xbar_demux_016:src0_channel -> tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_demux_016_src1_endofpacket                                                                   : std_logic;                      -- rsp_xbar_demux_016:src1_endofpacket -> cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_demux_016_src1_valid                                                                         : std_logic;                      -- rsp_xbar_demux_016:src1_valid -> cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_demux_016_src1_startofpacket                                                                 : std_logic;                      -- rsp_xbar_demux_016:src1_startofpacket -> cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_demux_016_src1_data                                                                          : std_logic_vector(96 downto 0);  -- rsp_xbar_demux_016:src1_data -> cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_demux_016_src1_channel                                                                       : std_logic_vector(1 downto 0);   -- rsp_xbar_demux_016:src1_channel -> cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:rp_channel
	signal addr_router_011_src_endofpacket                                                                       : std_logic;                      -- addr_router_011:src_endofpacket -> cmd_xbar_demux_011:sink_endofpacket
	signal addr_router_011_src_valid                                                                             : std_logic;                      -- addr_router_011:src_valid -> cmd_xbar_demux_011:sink_valid
	signal addr_router_011_src_startofpacket                                                                     : std_logic;                      -- addr_router_011:src_startofpacket -> cmd_xbar_demux_011:sink_startofpacket
	signal addr_router_011_src_data                                                                              : std_logic_vector(96 downto 0);  -- addr_router_011:src_data -> cmd_xbar_demux_011:sink_data
	signal addr_router_011_src_channel                                                                           : std_logic_vector(1 downto 0);   -- addr_router_011:src_channel -> cmd_xbar_demux_011:sink_channel
	signal addr_router_011_src_ready                                                                             : std_logic;                      -- cmd_xbar_demux_011:sink_ready -> addr_router_011:src_ready
	signal rsp_xbar_demux_016_src0_ready                                                                         : std_logic;                      -- tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_016:src0_ready
	signal addr_router_012_src_endofpacket                                                                       : std_logic;                      -- addr_router_012:src_endofpacket -> cmd_xbar_demux_012:sink_endofpacket
	signal addr_router_012_src_valid                                                                             : std_logic;                      -- addr_router_012:src_valid -> cmd_xbar_demux_012:sink_valid
	signal addr_router_012_src_startofpacket                                                                     : std_logic;                      -- addr_router_012:src_startofpacket -> cmd_xbar_demux_012:sink_startofpacket
	signal addr_router_012_src_data                                                                              : std_logic_vector(96 downto 0);  -- addr_router_012:src_data -> cmd_xbar_demux_012:sink_data
	signal addr_router_012_src_channel                                                                           : std_logic_vector(1 downto 0);   -- addr_router_012:src_channel -> cmd_xbar_demux_012:sink_channel
	signal addr_router_012_src_ready                                                                             : std_logic;                      -- cmd_xbar_demux_012:sink_ready -> addr_router_012:src_ready
	signal rsp_xbar_demux_016_src1_ready                                                                         : std_logic;                      -- cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_016:src1_ready
	signal cmd_xbar_demux_008_src0_ready                                                                         : std_logic;                      -- width_adapter:in_ready -> cmd_xbar_demux_008:src0_ready
	signal width_adapter_src_endofpacket                                                                         : std_logic;                      -- width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	signal width_adapter_src_valid                                                                               : std_logic;                      -- width_adapter:out_valid -> burst_adapter:sink0_valid
	signal width_adapter_src_startofpacket                                                                       : std_logic;                      -- width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	signal width_adapter_src_data                                                                                : std_logic_vector(76 downto 0);  -- width_adapter:out_data -> burst_adapter:sink0_data
	signal width_adapter_src_ready                                                                               : std_logic;                      -- burst_adapter:sink0_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                             : std_logic_vector(1 downto 0);   -- width_adapter:out_channel -> burst_adapter:sink0_channel
	signal id_router_013_src_endofpacket                                                                         : std_logic;                      -- id_router_013:src_endofpacket -> width_adapter_001:in_endofpacket
	signal id_router_013_src_valid                                                                               : std_logic;                      -- id_router_013:src_valid -> width_adapter_001:in_valid
	signal id_router_013_src_startofpacket                                                                       : std_logic;                      -- id_router_013:src_startofpacket -> width_adapter_001:in_startofpacket
	signal id_router_013_src_data                                                                                : std_logic_vector(76 downto 0);  -- id_router_013:src_data -> width_adapter_001:in_data
	signal id_router_013_src_channel                                                                             : std_logic_vector(1 downto 0);   -- id_router_013:src_channel -> width_adapter_001:in_channel
	signal id_router_013_src_ready                                                                               : std_logic;                      -- width_adapter_001:in_ready -> id_router_013:src_ready
	signal width_adapter_001_src_endofpacket                                                                     : std_logic;                      -- width_adapter_001:out_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	signal width_adapter_001_src_valid                                                                           : std_logic;                      -- width_adapter_001:out_valid -> rsp_xbar_demux_013:sink_valid
	signal width_adapter_001_src_startofpacket                                                                   : std_logic;                      -- width_adapter_001:out_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	signal width_adapter_001_src_data                                                                            : std_logic_vector(94 downto 0);  -- width_adapter_001:out_data -> rsp_xbar_demux_013:sink_data
	signal width_adapter_001_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_013:sink_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                         : std_logic_vector(1 downto 0);   -- width_adapter_001:out_channel -> rsp_xbar_demux_013:sink_channel
	signal cmd_xbar_demux_008_src1_ready                                                                         : std_logic;                      -- width_adapter_002:in_ready -> cmd_xbar_demux_008:src1_ready
	signal width_adapter_002_src_endofpacket                                                                     : std_logic;                      -- width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	signal width_adapter_002_src_valid                                                                           : std_logic;                      -- width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	signal width_adapter_002_src_startofpacket                                                                   : std_logic;                      -- width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	signal width_adapter_002_src_data                                                                            : std_logic_vector(76 downto 0);  -- width_adapter_002:out_data -> burst_adapter_001:sink0_data
	signal width_adapter_002_src_ready                                                                           : std_logic;                      -- burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	signal width_adapter_002_src_channel                                                                         : std_logic_vector(1 downto 0);   -- width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	signal id_router_014_src_endofpacket                                                                         : std_logic;                      -- id_router_014:src_endofpacket -> width_adapter_003:in_endofpacket
	signal id_router_014_src_valid                                                                               : std_logic;                      -- id_router_014:src_valid -> width_adapter_003:in_valid
	signal id_router_014_src_startofpacket                                                                       : std_logic;                      -- id_router_014:src_startofpacket -> width_adapter_003:in_startofpacket
	signal id_router_014_src_data                                                                                : std_logic_vector(76 downto 0);  -- id_router_014:src_data -> width_adapter_003:in_data
	signal id_router_014_src_channel                                                                             : std_logic_vector(1 downto 0);   -- id_router_014:src_channel -> width_adapter_003:in_channel
	signal id_router_014_src_ready                                                                               : std_logic;                      -- width_adapter_003:in_ready -> id_router_014:src_ready
	signal width_adapter_003_src_endofpacket                                                                     : std_logic;                      -- width_adapter_003:out_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	signal width_adapter_003_src_valid                                                                           : std_logic;                      -- width_adapter_003:out_valid -> rsp_xbar_demux_014:sink_valid
	signal width_adapter_003_src_startofpacket                                                                   : std_logic;                      -- width_adapter_003:out_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	signal width_adapter_003_src_data                                                                            : std_logic_vector(94 downto 0);  -- width_adapter_003:out_data -> rsp_xbar_demux_014:sink_data
	signal width_adapter_003_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_014:sink_ready -> width_adapter_003:out_ready
	signal width_adapter_003_src_channel                                                                         : std_logic_vector(1 downto 0);   -- width_adapter_003:out_channel -> rsp_xbar_demux_014:sink_channel
	signal cmd_xbar_mux_016_src_endofpacket                                                                      : std_logic;                      -- cmd_xbar_mux_016:src_endofpacket -> width_adapter_004:in_endofpacket
	signal cmd_xbar_mux_016_src_valid                                                                            : std_logic;                      -- cmd_xbar_mux_016:src_valid -> width_adapter_004:in_valid
	signal cmd_xbar_mux_016_src_startofpacket                                                                    : std_logic;                      -- cmd_xbar_mux_016:src_startofpacket -> width_adapter_004:in_startofpacket
	signal cmd_xbar_mux_016_src_data                                                                             : std_logic_vector(96 downto 0);  -- cmd_xbar_mux_016:src_data -> width_adapter_004:in_data
	signal cmd_xbar_mux_016_src_channel                                                                          : std_logic_vector(1 downto 0);   -- cmd_xbar_mux_016:src_channel -> width_adapter_004:in_channel
	signal cmd_xbar_mux_016_src_ready                                                                            : std_logic;                      -- width_adapter_004:in_ready -> cmd_xbar_mux_016:src_ready
	signal width_adapter_004_src_endofpacket                                                                     : std_logic;                      -- width_adapter_004:out_endofpacket -> sdram_0_avl_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal width_adapter_004_src_valid                                                                           : std_logic;                      -- width_adapter_004:out_valid -> sdram_0_avl_translator_avalon_universal_slave_0_agent:cp_valid
	signal width_adapter_004_src_startofpacket                                                                   : std_logic;                      -- width_adapter_004:out_startofpacket -> sdram_0_avl_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal width_adapter_004_src_data                                                                            : std_logic_vector(132 downto 0); -- width_adapter_004:out_data -> sdram_0_avl_translator_avalon_universal_slave_0_agent:cp_data
	signal width_adapter_004_src_ready                                                                           : std_logic;                      -- sdram_0_avl_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter_004:out_ready
	signal width_adapter_004_src_channel                                                                         : std_logic_vector(1 downto 0);   -- width_adapter_004:out_channel -> sdram_0_avl_translator_avalon_universal_slave_0_agent:cp_channel
	signal id_router_016_src_endofpacket                                                                         : std_logic;                      -- id_router_016:src_endofpacket -> width_adapter_005:in_endofpacket
	signal id_router_016_src_valid                                                                               : std_logic;                      -- id_router_016:src_valid -> width_adapter_005:in_valid
	signal id_router_016_src_startofpacket                                                                       : std_logic;                      -- id_router_016:src_startofpacket -> width_adapter_005:in_startofpacket
	signal id_router_016_src_data                                                                                : std_logic_vector(132 downto 0); -- id_router_016:src_data -> width_adapter_005:in_data
	signal id_router_016_src_channel                                                                             : std_logic_vector(1 downto 0);   -- id_router_016:src_channel -> width_adapter_005:in_channel
	signal id_router_016_src_ready                                                                               : std_logic;                      -- width_adapter_005:in_ready -> id_router_016:src_ready
	signal width_adapter_005_src_endofpacket                                                                     : std_logic;                      -- width_adapter_005:out_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	signal width_adapter_005_src_valid                                                                           : std_logic;                      -- width_adapter_005:out_valid -> rsp_xbar_demux_016:sink_valid
	signal width_adapter_005_src_startofpacket                                                                   : std_logic;                      -- width_adapter_005:out_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	signal width_adapter_005_src_data                                                                            : std_logic_vector(96 downto 0);  -- width_adapter_005:out_data -> rsp_xbar_demux_016:sink_data
	signal width_adapter_005_src_ready                                                                           : std_logic;                      -- rsp_xbar_demux_016:sink_ready -> width_adapter_005:out_ready
	signal width_adapter_005_src_channel                                                                         : std_logic_vector(1 downto 0);   -- width_adapter_005:out_channel -> rsp_xbar_demux_016:sink_channel
	signal limiter_cmd_valid_data                                                                                : std_logic_vector(3 downto 0);   -- limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	signal limiter_001_cmd_valid_data                                                                            : std_logic_vector(3 downto 0);   -- limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	signal limiter_002_cmd_valid_data                                                                            : std_logic_vector(7 downto 0);   -- limiter_002:cmd_src_valid -> cmd_xbar_demux_007:sink_valid
	signal limiter_003_cmd_valid_data                                                                            : std_logic_vector(1 downto 0);   -- limiter_003:cmd_src_valid -> cmd_xbar_demux_008:sink_valid
	signal linux_cpu_d_irq_irq                                                                                   : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> linux_cpu:d_irq
	signal irq_mapper_receiver0_irq                                                                              : std_logic;                      -- irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	signal irq_synchronizer_receiver_irq                                                                         : std_logic_vector(0 downto 0);   -- jtag_uart:av_irq -> irq_synchronizer:receiver_irq
	signal irq_mapper_receiver1_irq                                                                              : std_logic;                      -- irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	signal irq_synchronizer_001_receiver_irq                                                                     : std_logic_vector(0 downto 0);   -- sgdma_rx:csr_irq -> irq_synchronizer_001:receiver_irq
	signal irq_mapper_receiver2_irq                                                                              : std_logic;                      -- irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	signal irq_synchronizer_002_receiver_irq                                                                     : std_logic_vector(0 downto 0);   -- sgdma_tx:csr_irq -> irq_synchronizer_002:receiver_irq
	signal irq_mapper_receiver3_irq                                                                              : std_logic;                      -- irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	signal irq_synchronizer_003_receiver_irq                                                                     : std_logic_vector(0 downto 0);   -- linux_timer_1ms:irq -> irq_synchronizer_003:receiver_irq
	signal irq_mapper_receiver4_irq                                                                              : std_logic;                      -- irq_synchronizer_004:sender_irq -> irq_mapper:receiver4_irq
	signal irq_synchronizer_004_receiver_irq                                                                     : std_logic_vector(0 downto 0);   -- gtp_regif_0:irq -> irq_synchronizer_004:receiver_irq
	signal tse_mac_receive_endofpacket                                                                           : std_logic;                      -- tse_mac:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	signal tse_mac_receive_valid                                                                                 : std_logic;                      -- tse_mac:ff_rx_dval -> avalon_st_adapter:in_0_valid
	signal tse_mac_receive_startofpacket                                                                         : std_logic;                      -- tse_mac:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	signal tse_mac_receive_error                                                                                 : std_logic_vector(5 downto 0);   -- tse_mac:rx_err -> avalon_st_adapter:in_0_error
	signal tse_mac_receive_empty                                                                                 : std_logic_vector(1 downto 0);   -- tse_mac:ff_rx_mod -> avalon_st_adapter:in_0_empty
	signal tse_mac_receive_data                                                                                  : std_logic_vector(31 downto 0);  -- tse_mac:ff_rx_data -> avalon_st_adapter:in_0_data
	signal tse_mac_receive_ready                                                                                 : std_logic;                      -- avalon_st_adapter:in_0_ready -> tse_mac:ff_rx_rdy
	signal avalon_st_adapter_out_0_endofpacket                                                                   : std_logic;                      -- avalon_st_adapter:out_0_endofpacket -> sgdma_rx:in_endofpacket
	signal avalon_st_adapter_out_0_valid                                                                         : std_logic;                      -- avalon_st_adapter:out_0_valid -> sgdma_rx:in_valid
	signal avalon_st_adapter_out_0_startofpacket                                                                 : std_logic;                      -- avalon_st_adapter:out_0_startofpacket -> sgdma_rx:in_startofpacket
	signal avalon_st_adapter_out_0_error                                                                         : std_logic_vector(5 downto 0);   -- avalon_st_adapter:out_0_error -> sgdma_rx:in_error
	signal avalon_st_adapter_out_0_empty                                                                         : std_logic_vector(1 downto 0);   -- avalon_st_adapter:out_0_empty -> sgdma_rx:in_empty
	signal avalon_st_adapter_out_0_data                                                                          : std_logic_vector(31 downto 0);  -- avalon_st_adapter:out_0_data -> sgdma_rx:in_data
	signal avalon_st_adapter_out_0_ready                                                                         : std_logic;                      -- sgdma_rx:in_ready -> avalon_st_adapter:out_0_ready
	signal clk_in_reset_reset_n_ports_inv                                                                        : std_logic;                      -- clk_in_reset_reset_n:inv -> [rst_controller:reset_in2, rst_controller_001:reset_in2, rst_controller_002:reset_in0, rst_controller_003:reset_in1]
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                            : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> jtag_uart:av_write_n
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                             : std_logic;                      -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> jtag_uart:av_read_n
	signal linux_timer_1ms_s1_translator_avalon_anti_slave_0_write_ports_inv                                     : std_logic;                      -- linux_timer_1ms_s1_translator_avalon_anti_slave_0_write:inv -> linux_timer_1ms:write_n
	signal sdram_0_avl_translator_avalon_anti_slave_0_inv                                                        : std_logic;                      -- sdram_0_avl_waitrequest:inv -> sdram_0_avl_translator:av_waitrequest
	signal rst_controller_reset_out_reset_ports_inv                                                              : std_logic;                      -- rst_controller_reset_out_reset:inv -> [jtag_uart:rst_n, linux_timer_1ms:reset_n, sgdma_rx:system_reset_n, sgdma_tx:system_reset_n, sysid:reset_n]
	signal sdram_0_afi_reset_reset_ports_inv                                                                     : std_logic;                      -- sdram_0_afi_reset_reset:inv -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_003:reset_in0, rst_controller_004:reset_in0]
	signal rst_controller_001_reset_out_reset_ports_inv                                                          : std_logic;                      -- rst_controller_001_reset_out_reset:inv -> linux_cpu:reset_n
	signal rst_controller_002_reset_out_reset_ports_inv                                                          : std_logic;                      -- rst_controller_002_reset_out_reset:inv -> sdram_0:soft_reset_n

begin

	linux_timer_1ms : component sopc_system_linux_timer_1ms
		port map (
			clk        => sdram_0_afi_half_clk_clk,                                          --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                          -- reset.reset_n
			address    => linux_timer_1ms_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => linux_timer_1ms_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => linux_timer_1ms_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => linux_timer_1ms_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => linux_timer_1ms_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_synchronizer_003_receiver_irq(0)                               --   irq.irq
		);

	jtag_uart : component sopc_system_jtag_uart
		port map (
			clk            => sdram_0_afi_half_clk_clk,                                                   --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                                   --             reset.reset_n
			av_chipselect  => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_synchronizer_receiver_irq(0)                                            --               irq.irq
		);

	sgdma_rx : component sopc_system_sgdma_rx
		port map (
			clk                           => sdram_0_afi_half_clk_clk,                               --              clk.clk
			system_reset_n                => rst_controller_reset_out_reset_ports_inv,               --            reset.reset_n
			csr_chipselect                => sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect, --              csr.chipselect
			csr_address                   => sgdma_rx_csr_translator_avalon_anti_slave_0_address,    --                 .address
			csr_read                      => sgdma_rx_csr_translator_avalon_anti_slave_0_read,       --                 .read
			csr_write                     => sgdma_rx_csr_translator_avalon_anti_slave_0_write,      --                 .write
			csr_writedata                 => sgdma_rx_csr_translator_avalon_anti_slave_0_writedata,  --                 .writedata
			csr_readdata                  => sgdma_rx_csr_translator_avalon_anti_slave_0_readdata,   --                 .readdata
			descriptor_read_readdata      => sgdma_rx_descriptor_read_readdata,                      --  descriptor_read.readdata
			descriptor_read_readdatavalid => sgdma_rx_descriptor_read_readdatavalid,                 --                 .readdatavalid
			descriptor_read_waitrequest   => sgdma_rx_descriptor_read_waitrequest,                   --                 .waitrequest
			descriptor_read_address       => sgdma_rx_descriptor_read_address,                       --                 .address
			descriptor_read_read          => sgdma_rx_descriptor_read_read,                          --                 .read
			descriptor_write_waitrequest  => sgdma_rx_descriptor_write_waitrequest,                  -- descriptor_write.waitrequest
			descriptor_write_address      => sgdma_rx_descriptor_write_address,                      --                 .address
			descriptor_write_write        => sgdma_rx_descriptor_write_write,                        --                 .write
			descriptor_write_writedata    => sgdma_rx_descriptor_write_writedata,                    --                 .writedata
			csr_irq                       => irq_synchronizer_001_receiver_irq(0),                   --          csr_irq.irq
			in_startofpacket              => avalon_st_adapter_out_0_startofpacket,                  --               in.startofpacket
			in_endofpacket                => avalon_st_adapter_out_0_endofpacket,                    --                 .endofpacket
			in_data                       => avalon_st_adapter_out_0_data,                           --                 .data
			in_valid                      => avalon_st_adapter_out_0_valid,                          --                 .valid
			in_ready                      => avalon_st_adapter_out_0_ready,                          --                 .ready
			in_empty                      => avalon_st_adapter_out_0_empty,                          --                 .empty
			in_error                      => avalon_st_adapter_out_0_error,                          --                 .error
			m_write_waitrequest           => sgdma_rx_m_write_waitrequest,                           --          m_write.waitrequest
			m_write_address               => sgdma_rx_m_write_address,                               --                 .address
			m_write_write                 => sgdma_rx_m_write_write,                                 --                 .write
			m_write_writedata             => sgdma_rx_m_write_writedata,                             --                 .writedata
			m_write_byteenable            => sgdma_rx_m_write_byteenable                             --                 .byteenable
		);

	sgdma_tx : component sopc_system_sgdma_tx
		port map (
			clk                           => sdram_0_afi_half_clk_clk,                               --              clk.clk
			system_reset_n                => rst_controller_reset_out_reset_ports_inv,               --            reset.reset_n
			csr_chipselect                => sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect, --              csr.chipselect
			csr_address                   => sgdma_tx_csr_translator_avalon_anti_slave_0_address,    --                 .address
			csr_read                      => sgdma_tx_csr_translator_avalon_anti_slave_0_read,       --                 .read
			csr_write                     => sgdma_tx_csr_translator_avalon_anti_slave_0_write,      --                 .write
			csr_writedata                 => sgdma_tx_csr_translator_avalon_anti_slave_0_writedata,  --                 .writedata
			csr_readdata                  => sgdma_tx_csr_translator_avalon_anti_slave_0_readdata,   --                 .readdata
			descriptor_read_readdata      => sgdma_tx_descriptor_read_readdata,                      --  descriptor_read.readdata
			descriptor_read_readdatavalid => sgdma_tx_descriptor_read_readdatavalid,                 --                 .readdatavalid
			descriptor_read_waitrequest   => sgdma_tx_descriptor_read_waitrequest,                   --                 .waitrequest
			descriptor_read_address       => sgdma_tx_descriptor_read_address,                       --                 .address
			descriptor_read_read          => sgdma_tx_descriptor_read_read,                          --                 .read
			descriptor_write_waitrequest  => sgdma_tx_descriptor_write_waitrequest,                  -- descriptor_write.waitrequest
			descriptor_write_address      => sgdma_tx_descriptor_write_address,                      --                 .address
			descriptor_write_write        => sgdma_tx_descriptor_write_write,                        --                 .write
			descriptor_write_writedata    => sgdma_tx_descriptor_write_writedata,                    --                 .writedata
			csr_irq                       => irq_synchronizer_002_receiver_irq(0),                   --          csr_irq.irq
			m_read_readdata               => sgdma_tx_m_read_readdata,                               --           m_read.readdata
			m_read_readdatavalid          => sgdma_tx_m_read_readdatavalid,                          --                 .readdatavalid
			m_read_waitrequest            => sgdma_tx_m_read_waitrequest,                            --                 .waitrequest
			m_read_address                => sgdma_tx_m_read_address,                                --                 .address
			m_read_read                   => sgdma_tx_m_read_read,                                   --                 .read
			out_data                      => sgdma_tx_out_data,                                      --              out.data
			out_valid                     => sgdma_tx_out_valid,                                     --                 .valid
			out_ready                     => sgdma_tx_out_ready,                                     --                 .ready
			out_endofpacket               => sgdma_tx_out_endofpacket,                               --                 .endofpacket
			out_startofpacket             => sgdma_tx_out_startofpacket,                             --                 .startofpacket
			out_empty                     => sgdma_tx_out_empty,                                     --                 .empty
			out_error                     => sgdma_tx_out_error                                      --                 .error
		);

	descriptor_memory : component sopc_system_descriptor_memory
		port map (
			clk        => sdram_0_afi_half_clk_clk,                                       --   clk1.clk
			address    => descriptor_memory_s1_translator_avalon_anti_slave_0_address,    --     s1.address
			clken      => descriptor_memory_s1_translator_avalon_anti_slave_0_clken,      --       .clken
			chipselect => descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			write      => descriptor_memory_s1_translator_avalon_anti_slave_0_write,      --       .write
			readdata   => descriptor_memory_s1_translator_avalon_anti_slave_0_readdata,   --       .readdata
			writedata  => descriptor_memory_s1_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable => descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                                 -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                              --       .reset_req
		);

	linux_cpu : component sopc_system_linux_cpu
		port map (
			clk                                   => sdram_0_afi_clk_clk,                                                    --                                  clk.clk
			reset_n                               => rst_controller_001_reset_out_reset_ports_inv,                           --                              reset_n.reset_n
			d_address                             => linux_cpu_data_master_address,                                          --                          data_master.address
			d_byteenable                          => linux_cpu_data_master_byteenable,                                       --                                     .byteenable
			d_read                                => linux_cpu_data_master_read,                                             --                                     .read
			d_readdata                            => linux_cpu_data_master_readdata,                                         --                                     .readdata
			d_waitrequest                         => linux_cpu_data_master_waitrequest,                                      --                                     .waitrequest
			d_write                               => linux_cpu_data_master_write,                                            --                                     .write
			d_writedata                           => linux_cpu_data_master_writedata,                                        --                                     .writedata
			d_readdatavalid                       => linux_cpu_data_master_readdatavalid,                                    --                                     .readdatavalid
			jtag_debug_module_debugaccess_to_roms => linux_cpu_data_master_debugaccess,                                      --                                     .debugaccess
			i_address                             => linux_cpu_instruction_master_address,                                   --                   instruction_master.address
			i_read                                => linux_cpu_instruction_master_read,                                      --                                     .read
			i_readdata                            => linux_cpu_instruction_master_readdata,                                  --                                     .readdata
			i_waitrequest                         => linux_cpu_instruction_master_waitrequest,                               --                                     .waitrequest
			i_readdatavalid                       => linux_cpu_instruction_master_readdatavalid,                             --                                     .readdatavalid
			dcm0_readdata                         => linux_cpu_tightly_coupled_data_master_0_readdata,                       --        tightly_coupled_data_master_0.readdata
			dcm0_waitrequest                      => linux_cpu_tightly_coupled_data_master_0_waitrequest,                    --                                     .waitrequest
			dcm0_readdatavalid                    => linux_cpu_tightly_coupled_data_master_0_readdatavalid,                  --                                     .readdatavalid
			dcm0_address                          => linux_cpu_tightly_coupled_data_master_0_address,                        --                                     .address
			dcm0_read                             => linux_cpu_tightly_coupled_data_master_0_read,                           --                                     .read
			dcm0_clken                            => linux_cpu_tightly_coupled_data_master_0_clken,                          --                                     .clken
			dcm0_byteenable                       => linux_cpu_tightly_coupled_data_master_0_byteenable,                     --                                     .byteenable
			dcm0_write                            => linux_cpu_tightly_coupled_data_master_0_write,                          --                                     .write
			dcm0_writedata                        => linux_cpu_tightly_coupled_data_master_0_writedata,                      --                                     .writedata
			icm0_readdata                         => linux_cpu_tightly_coupled_instruction_master_0_readdata,                -- tightly_coupled_instruction_master_0.readdata
			icm0_waitrequest                      => linux_cpu_tightly_coupled_instruction_master_0_waitrequest,             --                                     .waitrequest
			icm0_readdatavalid                    => linux_cpu_tightly_coupled_instruction_master_0_readdatavalid,           --                                     .readdatavalid
			icm0_address                          => linux_cpu_tightly_coupled_instruction_master_0_address,                 --                                     .address
			icm0_read                             => linux_cpu_tightly_coupled_instruction_master_0_read,                    --                                     .read
			icm0_clken                            => linux_cpu_tightly_coupled_instruction_master_0_clken,                   --                                     .clken
			d_irq                                 => linux_cpu_d_irq_irq,                                                    --                                d_irq.irq
			jtag_debug_module_resetrequest        => linux_cpu_jtag_debug_module_reset_reset,                                --              jtag_debug_module_reset.reset
			jtag_debug_module_address             => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_address,     --                    jtag_debug_module.address
			jtag_debug_module_byteenable          => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,  --                                     .byteenable
			jtag_debug_module_debugaccess         => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess, --                                     .debugaccess
			jtag_debug_module_read                => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_read,        --                                     .read
			jtag_debug_module_readdata            => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata,    --                                     .readdata
			jtag_debug_module_waitrequest         => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest, --                                     .waitrequest
			jtag_debug_module_write               => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_write,       --                                     .write
			jtag_debug_module_writedata           => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata,   --                                     .writedata
			no_ci_readra                          => open                                                                    --            custom_instruction_master.readra
		);

	sysid : component sopc_system_sysid
		port map (
			clock    => sdram_0_afi_half_clk_clk,                                      --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                      --         reset.reset_n
			readdata => sysid_control_slave_translator_avalon_anti_slave_0_readdata,   -- control_slave.readdata
			address  => sysid_control_slave_translator_avalon_anti_slave_0_address(0)  --              .address
		);

	sdram_0 : component sopc_system_sdram_0
		port map (
			pll_ref_clk        => clk_in_clk,                                                    --      pll_ref_clk.clk
			global_reset_n     => clk_in_reset_reset_n,                                          --     global_reset.reset_n
			soft_reset_n       => rst_controller_002_reset_out_reset_ports_inv,                  --       soft_reset.reset_n
			afi_clk            => sdram_0_afi_clk_clk,                                           --          afi_clk.clk
			afi_half_clk       => sdram_0_afi_half_clk_clk,                                      --     afi_half_clk.clk
			afi_reset_n        => sdram_0_afi_reset_reset,                                       --        afi_reset.reset_n
			afi_reset_export_n => open,                                                          -- afi_reset_export.reset_n
			mem_a              => ddr2_mem_mem_a,                                                --           memory.mem_a
			mem_ba             => ddr2_mem_mem_ba,                                               --                 .mem_ba
			mem_ck             => ddr2_mem_mem_ck,                                               --                 .mem_ck
			mem_ck_n           => ddr2_mem_mem_ck_n,                                             --                 .mem_ck_n
			mem_cke            => ddr2_mem_mem_cke,                                              --                 .mem_cke
			mem_cs_n           => ddr2_mem_mem_cs_n,                                             --                 .mem_cs_n
			mem_dm             => ddr2_mem_mem_dm,                                               --                 .mem_dm
			mem_ras_n          => ddr2_mem_mem_ras_n,                                            --                 .mem_ras_n
			mem_cas_n          => ddr2_mem_mem_cas_n,                                            --                 .mem_cas_n
			mem_we_n           => ddr2_mem_mem_we_n,                                             --                 .mem_we_n
			mem_dq             => ddr2_mem_mem_dq,                                               --                 .mem_dq
			mem_dqs            => ddr2_mem_mem_dqs,                                              --                 .mem_dqs
			mem_dqs_n          => ddr2_mem_mem_dqs_n,                                            --                 .mem_dqs_n
			mem_odt            => ddr2_mem_mem_odt,                                              --                 .mem_odt
			avl_ready          => sdram_0_avl_waitrequest,                                       --              avl.waitrequest_n
			avl_burstbegin     => sdram_0_avl_translator_avalon_anti_slave_0_beginbursttransfer, --                 .beginbursttransfer
			avl_addr           => sdram_0_avl_translator_avalon_anti_slave_0_address,            --                 .address
			avl_rdata_valid    => sdram_0_avl_translator_avalon_anti_slave_0_readdatavalid,      --                 .readdatavalid
			avl_rdata          => sdram_0_avl_translator_avalon_anti_slave_0_readdata,           --                 .readdata
			avl_wdata          => sdram_0_avl_translator_avalon_anti_slave_0_writedata,          --                 .writedata
			avl_be             => sdram_0_avl_translator_avalon_anti_slave_0_byteenable,         --                 .byteenable
			avl_read_req       => sdram_0_avl_translator_avalon_anti_slave_0_read,               --                 .read
			avl_write_req      => sdram_0_avl_translator_avalon_anti_slave_0_write,              --                 .write
			avl_size           => sdram_0_avl_translator_avalon_anti_slave_0_burstcount,         --                 .burstcount
			local_init_done    => ddr2_status_local_init_done,                                   --           status.local_init_done
			local_cal_success  => ddr2_status_local_cal_success,                                 --                 .local_cal_success
			local_cal_fail     => ddr2_status_local_cal_fail,                                    --                 .local_cal_fail
			oct_rdn            => ddr2_oct_rdn,                                                  --              oct.rdn
			oct_rup            => ddr2_oct_rup                                                   --                 .rup
		);

	cfi_flash_ts_controller : component sopc_system_cfi_flash_ts_controller
		generic map (
			TCM_ADDRESS_W                  => 27,
			TCM_DATA_W                     => 16,
			TCM_BYTEENABLE_W               => 2,
			TCM_READ_WAIT                  => 230,
			TCM_WRITE_WAIT                 => 230,
			TCM_SETUP_WAIT                 => 65,
			TCM_DATA_HOLD                  => 35,
			TCM_TURNAROUND_TIME            => 2,
			TCM_TIMING_UNITS               => 0,
			TCM_READLATENCY                => 2,
			TCM_SYMBOLS_PER_WORD           => 2,
			USE_READDATA                   => 1,
			USE_WRITEDATA                  => 1,
			USE_READ                       => 0,
			USE_WRITE                      => 1,
			USE_BYTEENABLE                 => 0,
			USE_CHIPSELECT                 => 1,
			USE_LOCK                       => 0,
			USE_ADDRESS                    => 1,
			USE_WAITREQUEST                => 0,
			USE_WRITEBYTEENABLE            => 0,
			USE_OUTPUTENABLE               => 1,
			USE_RESETREQUEST               => 0,
			USE_IRQ                        => 0,
			USE_RESET_OUTPUT               => 1,
			ACTIVE_LOW_READ                => 1,
			ACTIVE_LOW_LOCK                => 0,
			ACTIVE_LOW_WRITE               => 1,
			ACTIVE_LOW_CHIPSELECT          => 1,
			ACTIVE_LOW_BYTEENABLE          => 0,
			ACTIVE_LOW_OUTPUTENABLE        => 1,
			ACTIVE_LOW_WRITEBYTEENABLE     => 0,
			ACTIVE_LOW_WAITREQUEST         => 0,
			ACTIVE_LOW_BEGINTRANSFER       => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0
		)
		port map (
			clk_clk                => sdram_0_afi_half_clk_clk,                                                 --   clk.clk
			reset_reset            => rst_controller_reset_out_reset,                                           -- reset.reset
			uas_address            => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_address,       --   uas.address
			uas_burstcount         => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_burstcount,    --      .burstcount
			uas_read               => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_read,          --      .read
			uas_write              => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_write,         --      .write
			uas_waitrequest        => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_waitrequest,   --      .waitrequest
			uas_readdatavalid      => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_readdatavalid, --      .readdatavalid
			uas_byteenable         => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_byteenable,    --      .byteenable
			uas_readdata           => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_readdata,      --      .readdata
			uas_writedata          => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_writedata,     --      .writedata
			uas_lock               => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_lock,          --      .lock
			uas_debugaccess        => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_debugaccess,   --      .debugaccess
			tcm_write_n_out        => cfi_flash_ts_controller_tcm_write_n_out,                                  --   tcm.write_n_out
			tcm_chipselect_n_out   => cfi_flash_ts_controller_tcm_chipselect_n_out,                             --      .chipselect_n_out
			tcm_outputenable_n_out => cfi_flash_ts_controller_tcm_outputenable_n_out,                           --      .outputenable_n_out
			tcm_reset_n_out        => cfi_flash_ts_controller_tcm_reset_n_out,                                  --      .reset_n_out
			tcm_request            => cfi_flash_ts_controller_tcm_request,                                      --      .request
			tcm_grant              => cfi_flash_ts_controller_tcm_grant,                                        --      .grant
			tcm_address_out        => cfi_flash_ts_controller_tcm_address_out,                                  --      .address_out
			tcm_data_out           => cfi_flash_ts_controller_tcm_data_out,                                     --      .data_out
			tcm_data_outen         => cfi_flash_ts_controller_tcm_data_outen,                                   --      .data_outen
			tcm_data_in            => cfi_flash_ts_controller_tcm_data_in                                       --      .data_in
		);

	cfi_flash_ts_bridge : component sopc_system_cfi_flash_ts_bridge
		port map (
			clk                           => sdram_0_afi_half_clk_clk,                       --   clk.clk
			reset                         => rst_controller_reset_out_reset,                 -- reset.reset
			request                       => cfi_flash_ts_controller_tcm_request,            --   tcs.request
			grant                         => cfi_flash_ts_controller_tcm_grant,              --      .grant
			tcs_tcm_address_out           => cfi_flash_ts_controller_tcm_address_out,        --      .address_out
			tcs_tcm_outputenable_n_out(0) => cfi_flash_ts_controller_tcm_outputenable_n_out, --      .outputenable_n_out
			tcs_tcm_reset_n_out(0)        => cfi_flash_ts_controller_tcm_reset_n_out,        --      .reset_n_out
			tcs_tcm_write_n_out(0)        => cfi_flash_ts_controller_tcm_write_n_out,        --      .write_n_out
			tcs_tcm_data_out              => cfi_flash_ts_controller_tcm_data_out,           --      .data_out
			tcs_tcm_data_outen            => cfi_flash_ts_controller_tcm_data_outen,         --      .data_outen
			tcs_tcm_data_in               => cfi_flash_ts_controller_tcm_data_in,            --      .data_in
			tcs_tcm_chipselect_n_out(0)   => cfi_flash_ts_controller_tcm_chipselect_n_out,   --      .chipselect_n_out
			tcm_address_out               => cfi_tcm_address_out,                            --   out.tcm_address_out
			tcm_outputenable_n_out        => cfi_tcm_outputenable_n_out,                     --      .tcm_outputenable_n_out
			tcm_reset_n_out               => cfi_tcm_reset_n_out,                            --      .tcm_reset_n_out
			tcm_write_n_out               => cfi_tcm_write_n_out,                            --      .tcm_write_n_out
			tcm_data_out                  => cfi_tcm_data_out,                               --      .tcm_data_out
			tcm_chipselect_n_out          => cfi_tcm_chipselect_n_out                        --      .tcm_chipselect_n_out
		);

	dma_to_descriptor_mem : component sopc_system_dma_to_descriptor_mem
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			ADDRESS_WIDTH     => 14,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => sdram_0_afi_half_clk_clk,                                              --   clk.clk
			reset            => rst_controller_reset_out_reset,                                        -- reset.reset
			s0_waitrequest   => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_waitrequest,   --    s0.waitrequest
			s0_readdata      => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_readdata,      --      .readdata
			s0_readdatavalid => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_readdatavalid, --      .readdatavalid
			s0_burstcount    => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_burstcount,    --      .burstcount
			s0_writedata     => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_writedata,     --      .writedata
			s0_address       => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_address,       --      .address
			s0_write         => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_write,         --      .write
			s0_read          => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_read,          --      .read
			s0_byteenable    => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_byteenable,    --      .byteenable
			s0_debugaccess   => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_debugaccess,   --      .debugaccess
			m0_waitrequest   => dma_to_descriptor_mem_m0_waitrequest,                                  --    m0.waitrequest
			m0_readdata      => dma_to_descriptor_mem_m0_readdata,                                     --      .readdata
			m0_readdatavalid => dma_to_descriptor_mem_m0_readdatavalid,                                --      .readdatavalid
			m0_burstcount    => dma_to_descriptor_mem_m0_burstcount,                                   --      .burstcount
			m0_writedata     => dma_to_descriptor_mem_m0_writedata,                                    --      .writedata
			m0_address       => dma_to_descriptor_mem_m0_address,                                      --      .address
			m0_write         => dma_to_descriptor_mem_m0_write,                                        --      .write
			m0_read          => dma_to_descriptor_mem_m0_read,                                         --      .read
			m0_byteenable    => dma_to_descriptor_mem_m0_byteenable,                                   --      .byteenable
			m0_debugaccess   => dma_to_descriptor_mem_m0_debugaccess                                   --      .debugaccess
		);

	gtp_regif_0 : component gtp_regif
		port map (
			avs_s0_address     => gtp_regif_0_s0_translator_avalon_anti_slave_0_address,     --               s0.address
			avs_s0_read        => gtp_regif_0_s0_translator_avalon_anti_slave_0_read,        --                 .read
			avs_s0_readdata    => gtp_regif_0_s0_translator_avalon_anti_slave_0_readdata,    --                 .readdata
			avs_s0_write       => gtp_regif_0_s0_translator_avalon_anti_slave_0_write,       --                 .write
			avs_s0_writedata   => gtp_regif_0_s0_translator_avalon_anti_slave_0_writedata,   --                 .writedata
			avs_s0_waitrequest => gtp_regif_0_s0_translator_avalon_anti_slave_0_waitrequest, --                 .waitrequest
			clk                => sdram_0_afi_half_clk_clk,                                  --            clock.clk
			reset              => rst_controller_003_reset_out_reset,                        --            reset.reset
			BUS_CLK            => gtpbus_CLK,                                                --   conduit_gtpbus.export
			BUS_RESET          => gtpbus_RESET,                                              --                 .export
			BUS_DIN            => gtpbus_DIN,                                                --                 .export
			BUS_DOUT           => gtpbus_DOUT,                                               --                 .export
			BUS_WR             => gtpbus_WR,                                                 --                 .export
			BUS_RD             => gtpbus_RD,                                                 --                 .export
			BUS_ACK            => gtpbus_ACK,                                                --                 .export
			BUS_ADDR           => gtpbus_ADDR,                                               --                 .export
			BUS_IRQ            => gtpbus_IRQ,                                                --                 .export
			irq                => irq_synchronizer_004_receiver_irq(0)                       -- interrupt_sender.irq
		);

	tse_mac : component sopc_system_tse_mac
		port map (
			clk           => sdram_0_afi_half_clk_clk,                                        -- control_port_clock_connection.clk
			reset         => rst_controller_reset_out_reset,                                  --              reset_connection.reset
			address       => tse_mac_control_port_translator_avalon_anti_slave_0_address,     --                  control_port.address
			readdata      => tse_mac_control_port_translator_avalon_anti_slave_0_readdata,    --                              .readdata
			read          => tse_mac_control_port_translator_avalon_anti_slave_0_read,        --                              .read
			writedata     => tse_mac_control_port_translator_avalon_anti_slave_0_writedata,   --                              .writedata
			write         => tse_mac_control_port_translator_avalon_anti_slave_0_write,       --                              .write
			waitrequest   => tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest, --                              .waitrequest
			tx_clk        => tse_txclk_clk,                                                   --   pcs_mac_tx_clock_connection.clk
			rx_clk        => tse_rxclk_clk,                                                   --   pcs_mac_rx_clock_connection.clk
			set_10        => tse_status_set_10,                                               --         mac_status_connection.set_10
			set_1000      => tse_status_set_1000,                                             --                              .set_1000
			eth_mode      => tse_status_eth_mode,                                             --                              .eth_mode
			ena_10        => tse_status_ena_10,                                               --                              .ena_10
			rgmii_in      => tse_rgmii_rgmii_in,                                              --          mac_rgmii_connection.rgmii_in
			rgmii_out     => tse_rgmii_rgmii_out,                                             --                              .rgmii_out
			rx_control    => tse_rgmii_rx_control,                                            --                              .rx_control
			tx_control    => tse_rgmii_tx_control,                                            --                              .tx_control
			ff_rx_clk     => sdram_0_afi_half_clk_clk,                                        --     transmit_clock_connection.clk
			ff_tx_clk     => sdram_0_afi_half_clk_clk,                                        --      receive_clock_connection.clk
			ff_rx_data    => tse_mac_receive_data,                                            --                       receive.data
			ff_rx_eop     => tse_mac_receive_endofpacket,                                     --                              .endofpacket
			rx_err        => tse_mac_receive_error,                                           --                              .error
			ff_rx_mod     => tse_mac_receive_empty,                                           --                              .empty
			ff_rx_rdy     => tse_mac_receive_ready,                                           --                              .ready
			ff_rx_sop     => tse_mac_receive_startofpacket,                                   --                              .startofpacket
			ff_rx_dval    => tse_mac_receive_valid,                                           --                              .valid
			ff_tx_data    => sgdma_tx_out_data,                                               --                      transmit.data
			ff_tx_eop     => sgdma_tx_out_endofpacket,                                        --                              .endofpacket
			ff_tx_err     => sgdma_tx_out_error,                                              --                              .error
			ff_tx_mod     => sgdma_tx_out_empty,                                              --                              .empty
			ff_tx_rdy     => sgdma_tx_out_ready,                                              --                              .ready
			ff_tx_sop     => sgdma_tx_out_startofpacket,                                      --                              .startofpacket
			ff_tx_wren    => sgdma_tx_out_valid,                                              --                              .valid
			mdc           => tse_mdio_mdc,                                                    --           mac_mdio_connection.mdc
			mdio_in       => tse_mdio_mdio_in,                                                --                              .mdio_in
			mdio_out      => tse_mdio_mdio_out,                                               --                              .mdio_out
			mdio_oen      => tse_mdio_mdio_oen,                                               --                              .mdio_oen
			xon_gen       => tse_misc_xon_gen,                                                --           mac_misc_connection.xon_gen
			xoff_gen      => tse_misc_xoff_gen,                                               --                              .xoff_gen
			magic_wakeup  => tse_misc_magic_wakeup,                                           --                              .magic_wakeup
			magic_sleep_n => tse_misc_magic_sleep_n,                                          --                              .magic_sleep_n
			ff_tx_crc_fwd => tse_misc_ff_tx_crc_fwd,                                          --                              .ff_tx_crc_fwd
			ff_tx_septy   => tse_misc_ff_tx_septy,                                            --                              .ff_tx_septy
			tx_ff_uflow   => tse_misc_tx_ff_uflow,                                            --                              .tx_ff_uflow
			ff_tx_a_full  => tse_misc_ff_tx_a_full,                                           --                              .ff_tx_a_full
			ff_tx_a_empty => tse_misc_ff_tx_a_empty,                                          --                              .ff_tx_a_empty
			rx_err_stat   => tse_misc_rx_err_stat,                                            --                              .rx_err_stat
			rx_frm_type   => tse_misc_rx_frm_type,                                            --                              .rx_frm_type
			ff_rx_dsav    => tse_misc_ff_rx_dsav,                                             --                              .ff_rx_dsav
			ff_rx_a_full  => tse_misc_ff_rx_a_full,                                           --                              .ff_rx_a_full
			ff_rx_a_empty => tse_misc_ff_rx_a_empty                                           --                              .ff_rx_a_empty
		);

	cfi_flash_ts_bridge_fpga : component sopc_system_cfi_flash_ts_bridge_fpga
		port map (
			clk                           => sdram_0_afi_half_clk_clk,                            --   clk.clk
			reset                         => rst_controller_reset_out_reset,                      -- reset.reset
			request                       => cfi_flash_ts_controller_fpga_tcm_request,            --   tcs.request
			grant                         => cfi_flash_ts_controller_fpga_tcm_grant,              --      .grant
			tcs_tcm_address_out           => cfi_flash_ts_controller_fpga_tcm_address_out,        --      .address_out
			tcs_tcm_outputenable_n_out(0) => cfi_flash_ts_controller_fpga_tcm_outputenable_n_out, --      .outputenable_n_out
			tcs_tcm_reset_n_out(0)        => cfi_flash_ts_controller_fpga_tcm_reset_n_out,        --      .reset_n_out
			tcs_tcm_write_n_out(0)        => cfi_flash_ts_controller_fpga_tcm_write_n_out,        --      .write_n_out
			tcs_tcm_data_out              => cfi_flash_ts_controller_fpga_tcm_data_out,           --      .data_out
			tcs_tcm_data_outen            => cfi_flash_ts_controller_fpga_tcm_data_outen,         --      .data_outen
			tcs_tcm_data_in               => cfi_flash_ts_controller_fpga_tcm_data_in,            --      .data_in
			tcs_tcm_chipselect_n_out(0)   => cfi_flash_ts_controller_fpga_tcm_chipselect_n_out,   --      .chipselect_n_out
			tcm_address_out               => cfi_fpga_tcm_address_out,                            --   out.tcm_address_out
			tcm_outputenable_n_out        => cfi_fpga_tcm_outputenable_n_out,                     --      .tcm_outputenable_n_out
			tcm_reset_n_out               => cfi_fpga_tcm_reset_n_out,                            --      .tcm_reset_n_out
			tcm_write_n_out               => cfi_fpga_tcm_write_n_out,                            --      .tcm_write_n_out
			tcm_data_out                  => cfi_fpga_tcm_data_out,                               --      .tcm_data_out
			tcm_chipselect_n_out          => cfi_fpga_tcm_chipselect_n_out                        --      .tcm_chipselect_n_out
		);

	cfi_flash_ts_controller_fpga : component sopc_system_cfi_flash_ts_controller
		generic map (
			TCM_ADDRESS_W                  => 27,
			TCM_DATA_W                     => 16,
			TCM_BYTEENABLE_W               => 2,
			TCM_READ_WAIT                  => 230,
			TCM_WRITE_WAIT                 => 230,
			TCM_SETUP_WAIT                 => 65,
			TCM_DATA_HOLD                  => 35,
			TCM_TURNAROUND_TIME            => 2,
			TCM_TIMING_UNITS               => 0,
			TCM_READLATENCY                => 2,
			TCM_SYMBOLS_PER_WORD           => 2,
			USE_READDATA                   => 1,
			USE_WRITEDATA                  => 1,
			USE_READ                       => 0,
			USE_WRITE                      => 1,
			USE_BYTEENABLE                 => 0,
			USE_CHIPSELECT                 => 1,
			USE_LOCK                       => 0,
			USE_ADDRESS                    => 1,
			USE_WAITREQUEST                => 0,
			USE_WRITEBYTEENABLE            => 0,
			USE_OUTPUTENABLE               => 1,
			USE_RESETREQUEST               => 0,
			USE_IRQ                        => 0,
			USE_RESET_OUTPUT               => 1,
			ACTIVE_LOW_READ                => 1,
			ACTIVE_LOW_LOCK                => 0,
			ACTIVE_LOW_WRITE               => 1,
			ACTIVE_LOW_CHIPSELECT          => 1,
			ACTIVE_LOW_BYTEENABLE          => 0,
			ACTIVE_LOW_OUTPUTENABLE        => 1,
			ACTIVE_LOW_WRITEBYTEENABLE     => 0,
			ACTIVE_LOW_WAITREQUEST         => 0,
			ACTIVE_LOW_BEGINTRANSFER       => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0
		)
		port map (
			clk_clk                => sdram_0_afi_half_clk_clk,                                                      --   clk.clk
			reset_reset            => rst_controller_reset_out_reset,                                                -- reset.reset
			uas_address            => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_address,       --   uas.address
			uas_burstcount         => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_burstcount,    --      .burstcount
			uas_read               => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_read,          --      .read
			uas_write              => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_write,         --      .write
			uas_waitrequest        => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_waitrequest,   --      .waitrequest
			uas_readdatavalid      => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_readdatavalid, --      .readdatavalid
			uas_byteenable         => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_byteenable,    --      .byteenable
			uas_readdata           => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_readdata,      --      .readdata
			uas_writedata          => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_writedata,     --      .writedata
			uas_lock               => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_lock,          --      .lock
			uas_debugaccess        => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_debugaccess,   --      .debugaccess
			tcm_write_n_out        => cfi_flash_ts_controller_fpga_tcm_write_n_out,                                  --   tcm.write_n_out
			tcm_chipselect_n_out   => cfi_flash_ts_controller_fpga_tcm_chipselect_n_out,                             --      .chipselect_n_out
			tcm_outputenable_n_out => cfi_flash_ts_controller_fpga_tcm_outputenable_n_out,                           --      .outputenable_n_out
			tcm_reset_n_out        => cfi_flash_ts_controller_fpga_tcm_reset_n_out,                                  --      .reset_n_out
			tcm_request            => cfi_flash_ts_controller_fpga_tcm_request,                                      --      .request
			tcm_grant              => cfi_flash_ts_controller_fpga_tcm_grant,                                        --      .grant
			tcm_address_out        => cfi_flash_ts_controller_fpga_tcm_address_out,                                  --      .address_out
			tcm_data_out           => cfi_flash_ts_controller_fpga_tcm_data_out,                                     --      .data_out
			tcm_data_outen         => cfi_flash_ts_controller_fpga_tcm_data_outen,                                   --      .data_outen
			tcm_data_in            => cfi_flash_ts_controller_fpga_tcm_data_in                                       --      .data_in
		);

	tse_dma_to_sdram_ccb : component sopc_system_tse_dma_to_sdram_ccb
		generic map (
			DATA_WIDTH          => 32,
			SYMBOL_WIDTH        => 8,
			ADDRESS_WIDTH       => 27,
			BURSTCOUNT_WIDTH    => 1,
			COMMAND_FIFO_DEPTH  => 4,
			RESPONSE_FIFO_DEPTH => 4,
			MASTER_SYNC_DEPTH   => 2,
			SLAVE_SYNC_DEPTH    => 2
		)
		port map (
			m0_clk           => sdram_0_afi_clk_clk,                                                  --   m0_clk.clk
			m0_reset         => rst_controller_001_reset_out_reset,                                   -- m0_reset.reset
			s0_clk           => sdram_0_afi_half_clk_clk,                                             --   s0_clk.clk
			s0_reset         => rst_controller_reset_out_reset,                                       -- s0_reset.reset
			s0_waitrequest   => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_waitrequest,   --       s0.waitrequest
			s0_readdata      => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_readdata,      --         .readdata
			s0_readdatavalid => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_readdatavalid, --         .readdatavalid
			s0_burstcount    => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_burstcount,    --         .burstcount
			s0_writedata     => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_writedata,     --         .writedata
			s0_address       => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_address,       --         .address
			s0_write         => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_write,         --         .write
			s0_read          => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_read,          --         .read
			s0_byteenable    => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_byteenable,    --         .byteenable
			s0_debugaccess   => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_debugaccess,   --         .debugaccess
			m0_waitrequest   => tse_dma_to_sdram_ccb_m0_waitrequest,                                  --       m0.waitrequest
			m0_readdata      => tse_dma_to_sdram_ccb_m0_readdata,                                     --         .readdata
			m0_readdatavalid => tse_dma_to_sdram_ccb_m0_readdatavalid,                                --         .readdatavalid
			m0_burstcount    => tse_dma_to_sdram_ccb_m0_burstcount,                                   --         .burstcount
			m0_writedata     => tse_dma_to_sdram_ccb_m0_writedata,                                    --         .writedata
			m0_address       => tse_dma_to_sdram_ccb_m0_address,                                      --         .address
			m0_write         => tse_dma_to_sdram_ccb_m0_write,                                        --         .write
			m0_read          => tse_dma_to_sdram_ccb_m0_read,                                         --         .read
			m0_byteenable    => tse_dma_to_sdram_ccb_m0_byteenable,                                   --         .byteenable
			m0_debugaccess   => tse_dma_to_sdram_ccb_m0_debugaccess                                   --         .debugaccess
		);

	cpu_to_peripherals_ccb : component sopc_system_cpu_to_peripherals_ccb
		generic map (
			DATA_WIDTH          => 32,
			SYMBOL_WIDTH        => 8,
			ADDRESS_WIDTH       => 23,
			BURSTCOUNT_WIDTH    => 1,
			COMMAND_FIFO_DEPTH  => 4,
			RESPONSE_FIFO_DEPTH => 4,
			MASTER_SYNC_DEPTH   => 2,
			SLAVE_SYNC_DEPTH    => 2
		)
		port map (
			m0_clk           => sdram_0_afi_half_clk_clk,                                               --   m0_clk.clk
			m0_reset         => rst_controller_reset_out_reset,                                         -- m0_reset.reset
			s0_clk           => sdram_0_afi_clk_clk,                                                    --   s0_clk.clk
			s0_reset         => rst_controller_001_reset_out_reset,                                     -- s0_reset.reset
			s0_waitrequest   => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_waitrequest,   --       s0.waitrequest
			s0_readdata      => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_readdata,      --         .readdata
			s0_readdatavalid => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_readdatavalid, --         .readdatavalid
			s0_burstcount    => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_burstcount,    --         .burstcount
			s0_writedata     => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_writedata,     --         .writedata
			s0_address       => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_address,       --         .address
			s0_write         => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_write,         --         .write
			s0_read          => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_read,          --         .read
			s0_byteenable    => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_byteenable,    --         .byteenable
			s0_debugaccess   => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_debugaccess,   --         .debugaccess
			m0_waitrequest   => cpu_to_peripherals_ccb_m0_waitrequest,                                  --       m0.waitrequest
			m0_readdata      => cpu_to_peripherals_ccb_m0_readdata,                                     --         .readdata
			m0_readdatavalid => cpu_to_peripherals_ccb_m0_readdatavalid,                                --         .readdatavalid
			m0_burstcount    => cpu_to_peripherals_ccb_m0_burstcount,                                   --         .burstcount
			m0_writedata     => cpu_to_peripherals_ccb_m0_writedata,                                    --         .writedata
			m0_address       => cpu_to_peripherals_ccb_m0_address,                                      --         .address
			m0_write         => cpu_to_peripherals_ccb_m0_write,                                        --         .write
			m0_read          => cpu_to_peripherals_ccb_m0_read,                                         --         .read
			m0_byteenable    => cpu_to_peripherals_ccb_m0_byteenable,                                   --         .byteenable
			m0_debugaccess   => cpu_to_peripherals_ccb_m0_debugaccess                                   --         .debugaccess
		);

	cpu_to_flash_ccb : component sopc_system_cpu_to_flash_ccb
		generic map (
			DATA_WIDTH          => 32,
			SYMBOL_WIDTH        => 8,
			ADDRESS_WIDTH       => 28,
			BURSTCOUNT_WIDTH    => 1,
			COMMAND_FIFO_DEPTH  => 4,
			RESPONSE_FIFO_DEPTH => 4,
			MASTER_SYNC_DEPTH   => 2,
			SLAVE_SYNC_DEPTH    => 2
		)
		port map (
			m0_clk           => sdram_0_afi_half_clk_clk,                                         --   m0_clk.clk
			m0_reset         => rst_controller_reset_out_reset,                                   -- m0_reset.reset
			s0_clk           => sdram_0_afi_clk_clk,                                              --   s0_clk.clk
			s0_reset         => rst_controller_001_reset_out_reset,                               -- s0_reset.reset
			s0_waitrequest   => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_waitrequest,   --       s0.waitrequest
			s0_readdata      => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_readdata,      --         .readdata
			s0_readdatavalid => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_readdatavalid, --         .readdatavalid
			s0_burstcount    => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_burstcount,    --         .burstcount
			s0_writedata     => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_writedata,     --         .writedata
			s0_address       => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_address,       --         .address
			s0_write         => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_write,         --         .write
			s0_read          => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_read,          --         .read
			s0_byteenable    => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_byteenable,    --         .byteenable
			s0_debugaccess   => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_debugaccess,   --         .debugaccess
			m0_waitrequest   => cpu_to_flash_ccb_m0_waitrequest,                                  --       m0.waitrequest
			m0_readdata      => cpu_to_flash_ccb_m0_readdata,                                     --         .readdata
			m0_readdatavalid => cpu_to_flash_ccb_m0_readdatavalid,                                --         .readdatavalid
			m0_burstcount    => cpu_to_flash_ccb_m0_burstcount,                                   --         .burstcount
			m0_writedata     => cpu_to_flash_ccb_m0_writedata,                                    --         .writedata
			m0_address       => cpu_to_flash_ccb_m0_address,                                      --         .address
			m0_write         => cpu_to_flash_ccb_m0_write,                                        --         .write
			m0_read          => cpu_to_flash_ccb_m0_read,                                         --         .read
			m0_byteenable    => cpu_to_flash_ccb_m0_byteenable,                                   --         .byteenable
			m0_debugaccess   => cpu_to_flash_ccb_m0_debugaccess                                   --         .debugaccess
		);

	cpu_to_sdram_pb : component sopc_system_cpu_to_sdram_pb
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			ADDRESS_WIDTH     => 27,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => sdram_0_afi_clk_clk,                                             --   clk.clk
			reset            => rst_controller_001_reset_out_reset,                              -- reset.reset
			s0_waitrequest   => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_waitrequest,   --    s0.waitrequest
			s0_readdata      => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_readdata,      --      .readdata
			s0_readdatavalid => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_readdatavalid, --      .readdatavalid
			s0_burstcount    => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_burstcount,    --      .burstcount
			s0_writedata     => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_writedata,     --      .writedata
			s0_address       => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_address,       --      .address
			s0_write         => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_write,         --      .write
			s0_read          => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_read,          --      .read
			s0_byteenable    => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_byteenable,    --      .byteenable
			s0_debugaccess   => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_debugaccess,   --      .debugaccess
			m0_waitrequest   => cpu_to_sdram_pb_m0_waitrequest,                                  --    m0.waitrequest
			m0_readdata      => cpu_to_sdram_pb_m0_readdata,                                     --      .readdata
			m0_readdatavalid => cpu_to_sdram_pb_m0_readdatavalid,                                --      .readdatavalid
			m0_burstcount    => cpu_to_sdram_pb_m0_burstcount,                                   --      .burstcount
			m0_writedata     => cpu_to_sdram_pb_m0_writedata,                                    --      .writedata
			m0_address       => cpu_to_sdram_pb_m0_address,                                      --      .address
			m0_write         => cpu_to_sdram_pb_m0_write,                                        --      .write
			m0_read          => cpu_to_sdram_pb_m0_read,                                         --      .read
			m0_byteenable    => cpu_to_sdram_pb_m0_byteenable,                                   --      .byteenable
			m0_debugaccess   => cpu_to_sdram_pb_m0_debugaccess                                   --      .debugaccess
		);

	tlb_miss_ram_1k : component sopc_system_tlb_miss_ram_1k
		port map (
			clk         => sdram_0_afi_clk_clk,                                          --   clk1.clk
			address     => tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_address,    --     s1.address
			clken       => tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_clken,      --       .clken
			chipselect  => tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			write       => tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_write,      --       .write
			readdata    => tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_readdata,   --       .readdata
			writedata   => tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable  => tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			reset       => rst_controller_001_reset_out_reset,                           -- reset1.reset
			reset_req   => rst_controller_001_reset_out_reset_req,                       --       .reset_req
			address2    => tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_address,    --     s2.address
			chipselect2 => tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			clken2      => tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_clken,      --       .clken
			write2      => tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_write,      --       .write
			readdata2   => tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_readdata,   --       .readdata
			writedata2  => tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable2 => tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			clk2        => sdram_0_afi_clk_clk,                                          --   clk2.clk
			reset2      => rst_controller_001_reset_out_reset,                           -- reset2.reset
			reset_req2  => rst_controller_001_reset_out_reset_req                        --       .reset_req
		);

	linux_cpu_data_master_translator : component sopc_system_linux_cpu_data_master_translator
		generic map (
			AV_ADDRESS_W                => 29,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 29,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => sdram_0_afi_clk_clk,                                                      --                       clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                       --                     reset.reset
			uav_address              => linux_cpu_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => linux_cpu_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => linux_cpu_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => linux_cpu_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => linux_cpu_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => linux_cpu_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => linux_cpu_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => linux_cpu_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => linux_cpu_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => linux_cpu_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => linux_cpu_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => linux_cpu_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => linux_cpu_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => linux_cpu_data_master_byteenable,                                         --                          .byteenable
			av_read                  => linux_cpu_data_master_read,                                               --                          .read
			av_readdata              => linux_cpu_data_master_readdata,                                           --                          .readdata
			av_readdatavalid         => linux_cpu_data_master_readdatavalid,                                      --                          .readdatavalid
			av_write                 => linux_cpu_data_master_write,                                              --                          .write
			av_writedata             => linux_cpu_data_master_writedata,                                          --                          .writedata
			av_debugaccess           => linux_cpu_data_master_debugaccess,                                        --                          .debugaccess
			av_burstcount            => "1",                                                                      --               (terminated)
			av_beginbursttransfer    => '0',                                                                      --               (terminated)
			av_begintransfer         => '0',                                                                      --               (terminated)
			av_chipselect            => '0',                                                                      --               (terminated)
			av_lock                  => '0',                                                                      --               (terminated)
			uav_clken                => open,                                                                     --               (terminated)
			av_clken                 => '1',                                                                      --               (terminated)
			uav_response             => "00",                                                                     --               (terminated)
			av_response              => open,                                                                     --               (terminated)
			uav_writeresponserequest => open,                                                                     --               (terminated)
			uav_writeresponsevalid   => '0',                                                                      --               (terminated)
			av_writeresponserequest  => '0',                                                                      --               (terminated)
			av_writeresponsevalid    => open                                                                      --               (terminated)
		);

	linux_cpu_instruction_master_translator : component sopc_system_linux_cpu_instruction_master_translator
		generic map (
			AV_ADDRESS_W                => 29,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 29,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 1,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => sdram_0_afi_clk_clk,                                                             --                       clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                              --                     reset.reset
			uav_address              => linux_cpu_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => linux_cpu_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => linux_cpu_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => linux_cpu_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => linux_cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => linux_cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => linux_cpu_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => linux_cpu_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => linux_cpu_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => linux_cpu_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => linux_cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => linux_cpu_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => linux_cpu_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read                  => linux_cpu_instruction_master_read,                                               --                          .read
			av_readdata              => linux_cpu_instruction_master_readdata,                                           --                          .readdata
			av_readdatavalid         => linux_cpu_instruction_master_readdatavalid,                                      --                          .readdatavalid
			av_burstcount            => "1",                                                                             --               (terminated)
			av_byteenable            => "1111",                                                                          --               (terminated)
			av_beginbursttransfer    => '0',                                                                             --               (terminated)
			av_begintransfer         => '0',                                                                             --               (terminated)
			av_chipselect            => '0',                                                                             --               (terminated)
			av_write                 => '0',                                                                             --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                              --               (terminated)
			av_lock                  => '0',                                                                             --               (terminated)
			av_debugaccess           => '0',                                                                             --               (terminated)
			uav_clken                => open,                                                                            --               (terminated)
			av_clken                 => '1',                                                                             --               (terminated)
			uav_response             => "00",                                                                            --               (terminated)
			av_response              => open,                                                                            --               (terminated)
			uav_writeresponserequest => open,                                                                            --               (terminated)
			uav_writeresponsevalid   => '0',                                                                             --               (terminated)
			av_writeresponserequest  => '0',                                                                             --               (terminated)
			av_writeresponsevalid    => open                                                                             --               (terminated)
		);

	linux_cpu_jtag_debug_module_translator : component sopc_system_linux_cpu_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 29,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_clk_clk,                                                                    --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                     --                    reset.reset
			uav_address              => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => linux_cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                                   --              (terminated)
			av_burstcount            => open,                                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                                   --              (terminated)
			av_lock                  => open,                                                                                   --              (terminated)
			av_chipselect            => open,                                                                                   --              (terminated)
			av_clken                 => open,                                                                                   --              (terminated)
			uav_clken                => '0',                                                                                    --              (terminated)
			av_outputenable          => open,                                                                                   --              (terminated)
			uav_response             => open,                                                                                   --              (terminated)
			av_response              => "00",                                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                                     --              (terminated)
		);

	cpu_to_flash_ccb_s0_translator : component sopc_system_cpu_to_flash_ccb_s0_translator
		generic map (
			AV_ADDRESS_W                   => 28,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 29,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 1,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_clk_clk,                                                            --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                             --                    reset.reset
			uav_address              => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_burstcount            => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_burstcount,                  --                         .burstcount
			av_byteenable            => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => cpu_to_flash_ccb_s0_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                           --              (terminated)
			av_beginbursttransfer    => open,                                                                           --              (terminated)
			av_writebyteenable       => open,                                                                           --              (terminated)
			av_lock                  => open,                                                                           --              (terminated)
			av_chipselect            => open,                                                                           --              (terminated)
			av_clken                 => open,                                                                           --              (terminated)
			uav_clken                => '0',                                                                            --              (terminated)
			av_outputenable          => open,                                                                           --              (terminated)
			uav_response             => open,                                                                           --              (terminated)
			av_response              => "00",                                                                           --              (terminated)
			uav_writeresponserequest => '0',                                                                            --              (terminated)
			uav_writeresponsevalid   => open,                                                                           --              (terminated)
			av_writeresponserequest  => open,                                                                           --              (terminated)
			av_writeresponsevalid    => '0'                                                                             --              (terminated)
		);

	cpu_to_peripherals_ccb_s0_translator : component sopc_system_cpu_to_peripherals_ccb_s0_translator
		generic map (
			AV_ADDRESS_W                   => 23,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 29,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 1,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_clk_clk,                                                                  --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                   --                    reset.reset
			uav_address              => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_burstcount            => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_burstcount,                  --                         .burstcount
			av_byteenable            => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => cpu_to_peripherals_ccb_s0_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                                 --              (terminated)
			av_writebyteenable       => open,                                                                                 --              (terminated)
			av_lock                  => open,                                                                                 --              (terminated)
			av_chipselect            => open,                                                                                 --              (terminated)
			av_clken                 => open,                                                                                 --              (terminated)
			uav_clken                => '0',                                                                                  --              (terminated)
			av_outputenable          => open,                                                                                 --              (terminated)
			uav_response             => open,                                                                                 --              (terminated)
			av_response              => "00",                                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                                   --              (terminated)
		);

	cpu_to_sdram_pb_s0_translator : component sopc_system_cpu_to_sdram_pb_s0_translator
		generic map (
			AV_ADDRESS_W                   => 27,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 29,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 1,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_clk_clk,                                                           --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                            --                    reset.reset
			uav_address              => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_burstcount            => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_burstcount,                  --                         .burstcount
			av_byteenable            => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => cpu_to_sdram_pb_s0_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                          --              (terminated)
			av_beginbursttransfer    => open,                                                                          --              (terminated)
			av_writebyteenable       => open,                                                                          --              (terminated)
			av_lock                  => open,                                                                          --              (terminated)
			av_chipselect            => open,                                                                          --              (terminated)
			av_clken                 => open,                                                                          --              (terminated)
			uav_clken                => '0',                                                                           --              (terminated)
			av_outputenable          => open,                                                                          --              (terminated)
			uav_response             => open,                                                                          --              (terminated)
			av_response              => "00",                                                                          --              (terminated)
			uav_writeresponserequest => '0',                                                                           --              (terminated)
			uav_writeresponsevalid   => open,                                                                          --              (terminated)
			av_writeresponserequest  => open,                                                                          --              (terminated)
			av_writeresponsevalid    => '0'                                                                            --              (terminated)
		);

	sgdma_tx_descriptor_write_translator : component sopc_system_sgdma_tx_descriptor_write_translator
		generic map (
			AV_ADDRESS_W                => 32,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 0,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                     --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                               --                     reset.reset
			uav_address              => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => sgdma_tx_descriptor_write_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => sgdma_tx_descriptor_write_waitrequest,                                        --                          .waitrequest
			av_write                 => sgdma_tx_descriptor_write_write,                                              --                          .write
			av_writedata             => sgdma_tx_descriptor_write_writedata,                                          --                          .writedata
			av_burstcount            => "1",                                                                          --               (terminated)
			av_byteenable            => "1111",                                                                       --               (terminated)
			av_beginbursttransfer    => '0',                                                                          --               (terminated)
			av_begintransfer         => '0',                                                                          --               (terminated)
			av_chipselect            => '0',                                                                          --               (terminated)
			av_read                  => '0',                                                                          --               (terminated)
			av_readdata              => open,                                                                         --               (terminated)
			av_readdatavalid         => open,                                                                         --               (terminated)
			av_lock                  => '0',                                                                          --               (terminated)
			av_debugaccess           => '0',                                                                          --               (terminated)
			uav_clken                => open,                                                                         --               (terminated)
			av_clken                 => '1',                                                                          --               (terminated)
			uav_response             => "00",                                                                         --               (terminated)
			av_response              => open,                                                                         --               (terminated)
			uav_writeresponserequest => open,                                                                         --               (terminated)
			uav_writeresponsevalid   => '0',                                                                          --               (terminated)
			av_writeresponserequest  => '0',                                                                          --               (terminated)
			av_writeresponsevalid    => open                                                                          --               (terminated)
		);

	sgdma_rx_descriptor_write_translator : component sopc_system_sgdma_tx_descriptor_write_translator
		generic map (
			AV_ADDRESS_W                => 32,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 0,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                     --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                               --                     reset.reset
			uav_address              => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => sgdma_rx_descriptor_write_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => sgdma_rx_descriptor_write_waitrequest,                                        --                          .waitrequest
			av_write                 => sgdma_rx_descriptor_write_write,                                              --                          .write
			av_writedata             => sgdma_rx_descriptor_write_writedata,                                          --                          .writedata
			av_burstcount            => "1",                                                                          --               (terminated)
			av_byteenable            => "1111",                                                                       --               (terminated)
			av_beginbursttransfer    => '0',                                                                          --               (terminated)
			av_begintransfer         => '0',                                                                          --               (terminated)
			av_chipselect            => '0',                                                                          --               (terminated)
			av_read                  => '0',                                                                          --               (terminated)
			av_readdata              => open,                                                                         --               (terminated)
			av_readdatavalid         => open,                                                                         --               (terminated)
			av_lock                  => '0',                                                                          --               (terminated)
			av_debugaccess           => '0',                                                                          --               (terminated)
			uav_clken                => open,                                                                         --               (terminated)
			av_clken                 => '1',                                                                          --               (terminated)
			uav_response             => "00",                                                                         --               (terminated)
			av_response              => open,                                                                         --               (terminated)
			uav_writeresponserequest => open,                                                                         --               (terminated)
			uav_writeresponsevalid   => '0',                                                                          --               (terminated)
			av_writeresponserequest  => '0',                                                                          --               (terminated)
			av_writeresponsevalid    => open                                                                          --               (terminated)
		);

	sgdma_rx_descriptor_read_translator : component sopc_system_sgdma_rx_descriptor_read_translator
		generic map (
			AV_ADDRESS_W                => 32,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                    --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                     reset.reset
			uav_address              => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => sgdma_rx_descriptor_read_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => sgdma_rx_descriptor_read_waitrequest,                                        --                          .waitrequest
			av_read                  => sgdma_rx_descriptor_read_read,                                               --                          .read
			av_readdata              => sgdma_rx_descriptor_read_readdata,                                           --                          .readdata
			av_readdatavalid         => sgdma_rx_descriptor_read_readdatavalid,                                      --                          .readdatavalid
			av_burstcount            => "1",                                                                         --               (terminated)
			av_byteenable            => "1111",                                                                      --               (terminated)
			av_beginbursttransfer    => '0',                                                                         --               (terminated)
			av_begintransfer         => '0',                                                                         --               (terminated)
			av_chipselect            => '0',                                                                         --               (terminated)
			av_write                 => '0',                                                                         --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                          --               (terminated)
			av_lock                  => '0',                                                                         --               (terminated)
			av_debugaccess           => '0',                                                                         --               (terminated)
			uav_clken                => open,                                                                        --               (terminated)
			av_clken                 => '1',                                                                         --               (terminated)
			uav_response             => "00",                                                                        --               (terminated)
			av_response              => open,                                                                        --               (terminated)
			uav_writeresponserequest => open,                                                                        --               (terminated)
			uav_writeresponsevalid   => '0',                                                                         --               (terminated)
			av_writeresponserequest  => '0',                                                                         --               (terminated)
			av_writeresponsevalid    => open                                                                         --               (terminated)
		);

	sgdma_tx_descriptor_read_translator : component sopc_system_sgdma_rx_descriptor_read_translator
		generic map (
			AV_ADDRESS_W                => 32,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                    --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                     reset.reset
			uav_address              => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => sgdma_tx_descriptor_read_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => sgdma_tx_descriptor_read_waitrequest,                                        --                          .waitrequest
			av_read                  => sgdma_tx_descriptor_read_read,                                               --                          .read
			av_readdata              => sgdma_tx_descriptor_read_readdata,                                           --                          .readdata
			av_readdatavalid         => sgdma_tx_descriptor_read_readdatavalid,                                      --                          .readdatavalid
			av_burstcount            => "1",                                                                         --               (terminated)
			av_byteenable            => "1111",                                                                      --               (terminated)
			av_beginbursttransfer    => '0',                                                                         --               (terminated)
			av_begintransfer         => '0',                                                                         --               (terminated)
			av_chipselect            => '0',                                                                         --               (terminated)
			av_write                 => '0',                                                                         --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                          --               (terminated)
			av_lock                  => '0',                                                                         --               (terminated)
			av_debugaccess           => '0',                                                                         --               (terminated)
			uav_clken                => open,                                                                        --               (terminated)
			av_clken                 => '1',                                                                         --               (terminated)
			uav_response             => "00",                                                                        --               (terminated)
			av_response              => open,                                                                        --               (terminated)
			uav_writeresponserequest => open,                                                                        --               (terminated)
			uav_writeresponsevalid   => '0',                                                                         --               (terminated)
			av_writeresponserequest  => '0',                                                                         --               (terminated)
			av_writeresponsevalid    => open                                                                         --               (terminated)
		);

	dma_to_descriptor_mem_s0_translator : component sopc_system_dma_to_descriptor_mem_s0_translator
		generic map (
			AV_ADDRESS_W                   => 14,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 1,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                            --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                      --                    reset.reset
			uav_address              => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_burstcount            => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_burstcount,                  --                         .burstcount
			av_byteenable            => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => dma_to_descriptor_mem_s0_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                                --              (terminated)
			av_beginbursttransfer    => open,                                                                                --              (terminated)
			av_writebyteenable       => open,                                                                                --              (terminated)
			av_lock                  => open,                                                                                --              (terminated)
			av_chipselect            => open,                                                                                --              (terminated)
			av_clken                 => open,                                                                                --              (terminated)
			uav_clken                => '0',                                                                                 --              (terminated)
			av_outputenable          => open,                                                                                --              (terminated)
			uav_response             => open,                                                                                --              (terminated)
			av_response              => "00",                                                                                --              (terminated)
			uav_writeresponserequest => '0',                                                                                 --              (terminated)
			uav_writeresponsevalid   => open,                                                                                --              (terminated)
			av_writeresponserequest  => open,                                                                                --              (terminated)
			av_writeresponsevalid    => '0'                                                                                  --              (terminated)
		);

	dma_to_descriptor_mem_m0_translator : component sopc_system_dma_to_descriptor_mem_m0_translator
		generic map (
			AV_ADDRESS_W                => 14,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 23,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 1,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                    --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                              --                     reset.reset
			uav_address              => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => dma_to_descriptor_mem_m0_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => dma_to_descriptor_mem_m0_waitrequest,                                        --                          .waitrequest
			av_burstcount            => dma_to_descriptor_mem_m0_burstcount,                                         --                          .burstcount
			av_byteenable            => dma_to_descriptor_mem_m0_byteenable,                                         --                          .byteenable
			av_read                  => dma_to_descriptor_mem_m0_read,                                               --                          .read
			av_readdata              => dma_to_descriptor_mem_m0_readdata,                                           --                          .readdata
			av_readdatavalid         => dma_to_descriptor_mem_m0_readdatavalid,                                      --                          .readdatavalid
			av_write                 => dma_to_descriptor_mem_m0_write,                                              --                          .write
			av_writedata             => dma_to_descriptor_mem_m0_writedata,                                          --                          .writedata
			av_debugaccess           => dma_to_descriptor_mem_m0_debugaccess,                                        --                          .debugaccess
			av_beginbursttransfer    => '0',                                                                         --               (terminated)
			av_begintransfer         => '0',                                                                         --               (terminated)
			av_chipselect            => '0',                                                                         --               (terminated)
			av_lock                  => '0',                                                                         --               (terminated)
			uav_clken                => open,                                                                        --               (terminated)
			av_clken                 => '1',                                                                         --               (terminated)
			uav_response             => "00",                                                                        --               (terminated)
			av_response              => open,                                                                        --               (terminated)
			uav_writeresponserequest => open,                                                                        --               (terminated)
			uav_writeresponsevalid   => '0',                                                                         --               (terminated)
			av_writeresponserequest  => '0',                                                                         --               (terminated)
			av_writeresponsevalid    => open                                                                         --               (terminated)
		);

	cpu_to_peripherals_ccb_m0_translator : component sopc_system_cpu_to_peripherals_ccb_m0_translator
		generic map (
			AV_ADDRESS_W                => 23,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 23,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 1,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                     --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                               --                     reset.reset
			uav_address              => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_to_peripherals_ccb_m0_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_to_peripherals_ccb_m0_waitrequest,                                        --                          .waitrequest
			av_burstcount            => cpu_to_peripherals_ccb_m0_burstcount,                                         --                          .burstcount
			av_byteenable            => cpu_to_peripherals_ccb_m0_byteenable,                                         --                          .byteenable
			av_read                  => cpu_to_peripherals_ccb_m0_read,                                               --                          .read
			av_readdata              => cpu_to_peripherals_ccb_m0_readdata,                                           --                          .readdata
			av_readdatavalid         => cpu_to_peripherals_ccb_m0_readdatavalid,                                      --                          .readdatavalid
			av_write                 => cpu_to_peripherals_ccb_m0_write,                                              --                          .write
			av_writedata             => cpu_to_peripherals_ccb_m0_writedata,                                          --                          .writedata
			av_debugaccess           => cpu_to_peripherals_ccb_m0_debugaccess,                                        --                          .debugaccess
			av_beginbursttransfer    => '0',                                                                          --               (terminated)
			av_begintransfer         => '0',                                                                          --               (terminated)
			av_chipselect            => '0',                                                                          --               (terminated)
			av_lock                  => '0',                                                                          --               (terminated)
			uav_clken                => open,                                                                         --               (terminated)
			av_clken                 => '1',                                                                          --               (terminated)
			uav_response             => "00",                                                                         --               (terminated)
			av_response              => open,                                                                         --               (terminated)
			uav_writeresponserequest => open,                                                                         --               (terminated)
			uav_writeresponsevalid   => '0',                                                                          --               (terminated)
			av_writeresponserequest  => '0',                                                                          --               (terminated)
			av_writeresponsevalid    => open                                                                          --               (terminated)
		);

	descriptor_memory_s1_translator : component sopc_system_descriptor_memory_s1_translator
		generic map (
			AV_ADDRESS_W                   => 11,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 23,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                        --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                  --                    reset.reset
			uav_address              => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => descriptor_memory_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => descriptor_memory_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => descriptor_memory_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => descriptor_memory_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => descriptor_memory_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect            => descriptor_memory_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_clken                 => descriptor_memory_s1_translator_avalon_anti_slave_0_clken,                       --                         .clken
			av_read                  => open,                                                                            --              (terminated)
			av_begintransfer         => open,                                                                            --              (terminated)
			av_beginbursttransfer    => open,                                                                            --              (terminated)
			av_burstcount            => open,                                                                            --              (terminated)
			av_readdatavalid         => '0',                                                                             --              (terminated)
			av_waitrequest           => '0',                                                                             --              (terminated)
			av_writebyteenable       => open,                                                                            --              (terminated)
			av_lock                  => open,                                                                            --              (terminated)
			uav_clken                => '0',                                                                             --              (terminated)
			av_debugaccess           => open,                                                                            --              (terminated)
			av_outputenable          => open,                                                                            --              (terminated)
			uav_response             => open,                                                                            --              (terminated)
			av_response              => "00",                                                                            --              (terminated)
			uav_writeresponserequest => '0',                                                                             --              (terminated)
			uav_writeresponsevalid   => open,                                                                            --              (terminated)
			av_writeresponserequest  => open,                                                                            --              (terminated)
			av_writeresponsevalid    => '0'                                                                              --              (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator : component sopc_system_jtag_uart_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 23,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                         --                    reset.reset
			uav_address              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                                   --              (terminated)
			av_burstcount            => open,                                                                                   --              (terminated)
			av_byteenable            => open,                                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                                   --              (terminated)
			av_lock                  => open,                                                                                   --              (terminated)
			av_clken                 => open,                                                                                   --              (terminated)
			uav_clken                => '0',                                                                                    --              (terminated)
			av_debugaccess           => open,                                                                                   --              (terminated)
			av_outputenable          => open,                                                                                   --              (terminated)
			uav_response             => open,                                                                                   --              (terminated)
			av_response              => "00",                                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                                     --              (terminated)
		);

	tse_mac_control_port_translator : component sopc_system_tse_mac_control_port_translator
		generic map (
			AV_ADDRESS_W                   => 8,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 23,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 1,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                        --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                  --                    reset.reset
			uav_address              => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => tse_mac_control_port_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => tse_mac_control_port_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => tse_mac_control_port_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => tse_mac_control_port_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => tse_mac_control_port_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => tse_mac_control_port_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_begintransfer         => open,                                                                            --              (terminated)
			av_beginbursttransfer    => open,                                                                            --              (terminated)
			av_burstcount            => open,                                                                            --              (terminated)
			av_byteenable            => open,                                                                            --              (terminated)
			av_readdatavalid         => '0',                                                                             --              (terminated)
			av_writebyteenable       => open,                                                                            --              (terminated)
			av_lock                  => open,                                                                            --              (terminated)
			av_chipselect            => open,                                                                            --              (terminated)
			av_clken                 => open,                                                                            --              (terminated)
			uav_clken                => '0',                                                                             --              (terminated)
			av_debugaccess           => open,                                                                            --              (terminated)
			av_outputenable          => open,                                                                            --              (terminated)
			uav_response             => open,                                                                            --              (terminated)
			av_response              => "00",                                                                            --              (terminated)
			uav_writeresponserequest => '0',                                                                             --              (terminated)
			uav_writeresponsevalid   => open,                                                                            --              (terminated)
			av_writeresponserequest  => open,                                                                            --              (terminated)
			av_writeresponsevalid    => '0'                                                                              --              (terminated)
		);

	sysid_control_slave_translator : component sopc_system_sysid_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 23,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                       --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                 --                    reset.reset
			uav_address              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sysid_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => sysid_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                           --              (terminated)
			av_read                  => open,                                                                           --              (terminated)
			av_writedata             => open,                                                                           --              (terminated)
			av_begintransfer         => open,                                                                           --              (terminated)
			av_beginbursttransfer    => open,                                                                           --              (terminated)
			av_burstcount            => open,                                                                           --              (terminated)
			av_byteenable            => open,                                                                           --              (terminated)
			av_readdatavalid         => '0',                                                                            --              (terminated)
			av_waitrequest           => '0',                                                                            --              (terminated)
			av_writebyteenable       => open,                                                                           --              (terminated)
			av_lock                  => open,                                                                           --              (terminated)
			av_chipselect            => open,                                                                           --              (terminated)
			av_clken                 => open,                                                                           --              (terminated)
			uav_clken                => '0',                                                                            --              (terminated)
			av_debugaccess           => open,                                                                           --              (terminated)
			av_outputenable          => open,                                                                           --              (terminated)
			uav_response             => open,                                                                           --              (terminated)
			av_response              => "00",                                                                           --              (terminated)
			uav_writeresponserequest => '0',                                                                            --              (terminated)
			uav_writeresponsevalid   => open,                                                                           --              (terminated)
			av_writeresponserequest  => open,                                                                           --              (terminated)
			av_writeresponsevalid    => '0'                                                                             --              (terminated)
		);

	linux_timer_1ms_s1_translator : component sopc_system_linux_timer_1ms_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 23,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                      --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                --                    reset.reset
			uav_address              => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => linux_timer_1ms_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => linux_timer_1ms_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => linux_timer_1ms_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => linux_timer_1ms_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => linux_timer_1ms_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                          --              (terminated)
			av_begintransfer         => open,                                                                          --              (terminated)
			av_beginbursttransfer    => open,                                                                          --              (terminated)
			av_burstcount            => open,                                                                          --              (terminated)
			av_byteenable            => open,                                                                          --              (terminated)
			av_readdatavalid         => '0',                                                                           --              (terminated)
			av_waitrequest           => '0',                                                                           --              (terminated)
			av_writebyteenable       => open,                                                                          --              (terminated)
			av_lock                  => open,                                                                          --              (terminated)
			av_clken                 => open,                                                                          --              (terminated)
			uav_clken                => '0',                                                                           --              (terminated)
			av_debugaccess           => open,                                                                          --              (terminated)
			av_outputenable          => open,                                                                          --              (terminated)
			uav_response             => open,                                                                          --              (terminated)
			av_response              => "00",                                                                          --              (terminated)
			uav_writeresponserequest => '0',                                                                           --              (terminated)
			uav_writeresponsevalid   => open,                                                                          --              (terminated)
			av_writeresponserequest  => open,                                                                          --              (terminated)
			av_writeresponsevalid    => '0'                                                                            --              (terminated)
		);

	gtp_regif_0_s0_translator : component sopc_system_gtp_regif_0_s0_translator
		generic map (
			AV_ADDRESS_W                   => 14,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 23,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                            --                    reset.reset
			uav_address              => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => gtp_regif_0_s0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => gtp_regif_0_s0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => gtp_regif_0_s0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => gtp_regif_0_s0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => gtp_regif_0_s0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => gtp_regif_0_s0_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_begintransfer         => open,                                                                      --              (terminated)
			av_beginbursttransfer    => open,                                                                      --              (terminated)
			av_burstcount            => open,                                                                      --              (terminated)
			av_byteenable            => open,                                                                      --              (terminated)
			av_readdatavalid         => '0',                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                      --              (terminated)
			av_lock                  => open,                                                                      --              (terminated)
			av_chipselect            => open,                                                                      --              (terminated)
			av_clken                 => open,                                                                      --              (terminated)
			uav_clken                => '0',                                                                       --              (terminated)
			av_debugaccess           => open,                                                                      --              (terminated)
			av_outputenable          => open,                                                                      --              (terminated)
			uav_response             => open,                                                                      --              (terminated)
			av_response              => "00",                                                                      --              (terminated)
			uav_writeresponserequest => '0',                                                                       --              (terminated)
			uav_writeresponsevalid   => open,                                                                      --              (terminated)
			av_writeresponserequest  => open,                                                                      --              (terminated)
			av_writeresponsevalid    => '0'                                                                        --              (terminated)
		);

	sgdma_tx_csr_translator : component sopc_system_sgdma_tx_csr_translator
		generic map (
			AV_ADDRESS_W                   => 4,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 23,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                          --                    reset.reset
			uav_address              => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sgdma_tx_csr_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sgdma_tx_csr_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => sgdma_tx_csr_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => sgdma_tx_csr_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sgdma_tx_csr_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => sgdma_tx_csr_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                    --              (terminated)
			av_beginbursttransfer    => open,                                                                    --              (terminated)
			av_burstcount            => open,                                                                    --              (terminated)
			av_byteenable            => open,                                                                    --              (terminated)
			av_readdatavalid         => '0',                                                                     --              (terminated)
			av_waitrequest           => '0',                                                                     --              (terminated)
			av_writebyteenable       => open,                                                                    --              (terminated)
			av_lock                  => open,                                                                    --              (terminated)
			av_clken                 => open,                                                                    --              (terminated)
			uav_clken                => '0',                                                                     --              (terminated)
			av_debugaccess           => open,                                                                    --              (terminated)
			av_outputenable          => open,                                                                    --              (terminated)
			uav_response             => open,                                                                    --              (terminated)
			av_response              => "00",                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                      --              (terminated)
		);

	sgdma_rx_csr_translator : component sopc_system_sgdma_tx_csr_translator
		generic map (
			AV_ADDRESS_W                   => 4,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 23,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                          --                    reset.reset
			uav_address              => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sgdma_rx_csr_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sgdma_rx_csr_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => sgdma_rx_csr_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => sgdma_rx_csr_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sgdma_rx_csr_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => sgdma_rx_csr_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                    --              (terminated)
			av_beginbursttransfer    => open,                                                                    --              (terminated)
			av_burstcount            => open,                                                                    --              (terminated)
			av_byteenable            => open,                                                                    --              (terminated)
			av_readdatavalid         => '0',                                                                     --              (terminated)
			av_waitrequest           => '0',                                                                     --              (terminated)
			av_writebyteenable       => open,                                                                    --              (terminated)
			av_lock                  => open,                                                                    --              (terminated)
			av_clken                 => open,                                                                    --              (terminated)
			uav_clken                => '0',                                                                     --              (terminated)
			av_debugaccess           => open,                                                                    --              (terminated)
			av_outputenable          => open,                                                                    --              (terminated)
			uav_response             => open,                                                                    --              (terminated)
			av_response              => "00",                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                      --              (terminated)
		);

	cpu_to_flash_ccb_m0_translator : component sopc_system_cpu_to_flash_ccb_m0_translator
		generic map (
			AV_ADDRESS_W                => 28,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 28,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 1,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                               --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                         --                     reset.reset
			uav_address              => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_to_flash_ccb_m0_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_to_flash_ccb_m0_waitrequest,                                        --                          .waitrequest
			av_burstcount            => cpu_to_flash_ccb_m0_burstcount,                                         --                          .burstcount
			av_byteenable            => cpu_to_flash_ccb_m0_byteenable,                                         --                          .byteenable
			av_read                  => cpu_to_flash_ccb_m0_read,                                               --                          .read
			av_readdata              => cpu_to_flash_ccb_m0_readdata,                                           --                          .readdata
			av_readdatavalid         => cpu_to_flash_ccb_m0_readdatavalid,                                      --                          .readdatavalid
			av_write                 => cpu_to_flash_ccb_m0_write,                                              --                          .write
			av_writedata             => cpu_to_flash_ccb_m0_writedata,                                          --                          .writedata
			av_debugaccess           => cpu_to_flash_ccb_m0_debugaccess,                                        --                          .debugaccess
			av_beginbursttransfer    => '0',                                                                    --               (terminated)
			av_begintransfer         => '0',                                                                    --               (terminated)
			av_chipselect            => '0',                                                                    --               (terminated)
			av_lock                  => '0',                                                                    --               (terminated)
			uav_clken                => open,                                                                   --               (terminated)
			av_clken                 => '1',                                                                    --               (terminated)
			uav_response             => "00",                                                                   --               (terminated)
			av_response              => open,                                                                   --               (terminated)
			uav_writeresponserequest => open,                                                                   --               (terminated)
			uav_writeresponsevalid   => '0',                                                                    --               (terminated)
			av_writeresponserequest  => '0',                                                                    --               (terminated)
			av_writeresponsevalid    => open                                                                    --               (terminated)
		);

	cfi_flash_ts_controller_fpga_uas_translator : component sopc_system_cfi_flash_ts_controller_fpga_uas_translator
		generic map (
			AV_ADDRESS_W                   => 27,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 2,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 28,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 1,
			AV_BURSTCOUNT_SYMBOLS          => 1,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                                    --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                              --                    reset.reset
			uav_address              => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_burstcount            => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_burstcount,                  --                         .burstcount
			av_byteenable            => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_lock                  => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_lock,                        --                         .lock
			av_debugaccess           => cfi_flash_ts_controller_fpga_uas_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                                        --              (terminated)
			av_beginbursttransfer    => open,                                                                                        --              (terminated)
			av_writebyteenable       => open,                                                                                        --              (terminated)
			av_chipselect            => open,                                                                                        --              (terminated)
			av_clken                 => open,                                                                                        --              (terminated)
			uav_clken                => '0',                                                                                         --              (terminated)
			av_outputenable          => open,                                                                                        --              (terminated)
			uav_response             => open,                                                                                        --              (terminated)
			av_response              => "00",                                                                                        --              (terminated)
			uav_writeresponserequest => '0',                                                                                         --              (terminated)
			uav_writeresponsevalid   => open,                                                                                        --              (terminated)
			av_writeresponserequest  => open,                                                                                        --              (terminated)
			av_writeresponsevalid    => '0'                                                                                          --              (terminated)
		);

	cfi_flash_ts_controller_uas_translator : component sopc_system_cfi_flash_ts_controller_fpga_uas_translator
		generic map (
			AV_ADDRESS_W                   => 27,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 2,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 28,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 1,
			AV_BURSTCOUNT_SYMBOLS          => 1,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                               --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                         --                    reset.reset
			uav_address              => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_burstcount            => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_burstcount,                  --                         .burstcount
			av_byteenable            => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_lock                  => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_lock,                        --                         .lock
			av_debugaccess           => cfi_flash_ts_controller_uas_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                                   --              (terminated)
			av_chipselect            => open,                                                                                   --              (terminated)
			av_clken                 => open,                                                                                   --              (terminated)
			uav_clken                => '0',                                                                                    --              (terminated)
			av_outputenable          => open,                                                                                   --              (terminated)
			uav_response             => open,                                                                                   --              (terminated)
			av_response              => "00",                                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                                     --              (terminated)
		);

	sgdma_tx_m_read_translator : component sopc_system_sgdma_rx_descriptor_read_translator
		generic map (
			AV_ADDRESS_W                => 32,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                           --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                     --                     reset.reset
			uav_address              => sgdma_tx_m_read_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => sgdma_tx_m_read_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => sgdma_tx_m_read_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => sgdma_tx_m_read_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => sgdma_tx_m_read_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => sgdma_tx_m_read_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => sgdma_tx_m_read_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => sgdma_tx_m_read_waitrequest,                                        --                          .waitrequest
			av_read                  => sgdma_tx_m_read_read,                                               --                          .read
			av_readdata              => sgdma_tx_m_read_readdata,                                           --                          .readdata
			av_readdatavalid         => sgdma_tx_m_read_readdatavalid,                                      --                          .readdatavalid
			av_burstcount            => "1",                                                                --               (terminated)
			av_byteenable            => "1111",                                                             --               (terminated)
			av_beginbursttransfer    => '0',                                                                --               (terminated)
			av_begintransfer         => '0',                                                                --               (terminated)
			av_chipselect            => '0',                                                                --               (terminated)
			av_write                 => '0',                                                                --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                 --               (terminated)
			av_lock                  => '0',                                                                --               (terminated)
			av_debugaccess           => '0',                                                                --               (terminated)
			uav_clken                => open,                                                               --               (terminated)
			av_clken                 => '1',                                                                --               (terminated)
			uav_response             => "00",                                                               --               (terminated)
			av_response              => open,                                                               --               (terminated)
			uav_writeresponserequest => open,                                                               --               (terminated)
			uav_writeresponsevalid   => '0',                                                                --               (terminated)
			av_writeresponserequest  => '0',                                                                --               (terminated)
			av_writeresponsevalid    => open                                                                --               (terminated)
		);

	sgdma_rx_m_write_translator : component sopc_system_sgdma_rx_m_write_translator
		generic map (
			AV_ADDRESS_W                => 32,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 32,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 0,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                            --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                      --                     reset.reset
			uav_address              => sgdma_rx_m_write_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => sgdma_rx_m_write_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => sgdma_rx_m_write_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => sgdma_rx_m_write_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => sgdma_rx_m_write_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => sgdma_rx_m_write_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => sgdma_rx_m_write_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => sgdma_rx_m_write_waitrequest,                                        --                          .waitrequest
			av_byteenable            => sgdma_rx_m_write_byteenable,                                         --                          .byteenable
			av_write                 => sgdma_rx_m_write_write,                                              --                          .write
			av_writedata             => sgdma_rx_m_write_writedata,                                          --                          .writedata
			av_burstcount            => "1",                                                                 --               (terminated)
			av_beginbursttransfer    => '0',                                                                 --               (terminated)
			av_begintransfer         => '0',                                                                 --               (terminated)
			av_chipselect            => '0',                                                                 --               (terminated)
			av_read                  => '0',                                                                 --               (terminated)
			av_readdata              => open,                                                                --               (terminated)
			av_readdatavalid         => open,                                                                --               (terminated)
			av_lock                  => '0',                                                                 --               (terminated)
			av_debugaccess           => '0',                                                                 --               (terminated)
			uav_clken                => open,                                                                --               (terminated)
			av_clken                 => '1',                                                                 --               (terminated)
			uav_response             => "00",                                                                --               (terminated)
			av_response              => open,                                                                --               (terminated)
			uav_writeresponserequest => open,                                                                --               (terminated)
			uav_writeresponsevalid   => '0',                                                                 --               (terminated)
			av_writeresponserequest  => '0',                                                                 --               (terminated)
			av_writeresponsevalid    => open                                                                 --               (terminated)
		);

	tse_dma_to_sdram_ccb_s0_translator : component sopc_system_tse_dma_to_sdram_ccb_s0_translator
		generic map (
			AV_ADDRESS_W                   => 27,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 32,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 1,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_half_clk_clk,                                                           --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                     --                    reset.reset
			uav_address              => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_burstcount            => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_burstcount,                  --                         .burstcount
			av_byteenable            => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => tse_dma_to_sdram_ccb_s0_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                               --              (terminated)
			av_beginbursttransfer    => open,                                                                               --              (terminated)
			av_writebyteenable       => open,                                                                               --              (terminated)
			av_lock                  => open,                                                                               --              (terminated)
			av_chipselect            => open,                                                                               --              (terminated)
			av_clken                 => open,                                                                               --              (terminated)
			uav_clken                => '0',                                                                                --              (terminated)
			av_outputenable          => open,                                                                               --              (terminated)
			uav_response             => open,                                                                               --              (terminated)
			av_response              => "00",                                                                               --              (terminated)
			uav_writeresponserequest => '0',                                                                                --              (terminated)
			uav_writeresponsevalid   => open,                                                                               --              (terminated)
			av_writeresponserequest  => open,                                                                               --              (terminated)
			av_writeresponsevalid    => '0'                                                                                 --              (terminated)
		);

	tse_dma_to_sdram_ccb_m0_translator : component sopc_system_tse_dma_to_sdram_ccb_m0_translator
		generic map (
			AV_ADDRESS_W                => 27,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 27,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 1,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => sdram_0_afi_clk_clk,                                                        --                       clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                         --                     reset.reset
			uav_address              => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => tse_dma_to_sdram_ccb_m0_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => tse_dma_to_sdram_ccb_m0_waitrequest,                                        --                          .waitrequest
			av_burstcount            => tse_dma_to_sdram_ccb_m0_burstcount,                                         --                          .burstcount
			av_byteenable            => tse_dma_to_sdram_ccb_m0_byteenable,                                         --                          .byteenable
			av_read                  => tse_dma_to_sdram_ccb_m0_read,                                               --                          .read
			av_readdata              => tse_dma_to_sdram_ccb_m0_readdata,                                           --                          .readdata
			av_readdatavalid         => tse_dma_to_sdram_ccb_m0_readdatavalid,                                      --                          .readdatavalid
			av_write                 => tse_dma_to_sdram_ccb_m0_write,                                              --                          .write
			av_writedata             => tse_dma_to_sdram_ccb_m0_writedata,                                          --                          .writedata
			av_debugaccess           => tse_dma_to_sdram_ccb_m0_debugaccess,                                        --                          .debugaccess
			av_beginbursttransfer    => '0',                                                                        --               (terminated)
			av_begintransfer         => '0',                                                                        --               (terminated)
			av_chipselect            => '0',                                                                        --               (terminated)
			av_lock                  => '0',                                                                        --               (terminated)
			uav_clken                => open,                                                                       --               (terminated)
			av_clken                 => '1',                                                                        --               (terminated)
			uav_response             => "00",                                                                       --               (terminated)
			av_response              => open,                                                                       --               (terminated)
			uav_writeresponserequest => open,                                                                       --               (terminated)
			uav_writeresponsevalid   => '0',                                                                        --               (terminated)
			av_writeresponserequest  => '0',                                                                        --               (terminated)
			av_writeresponsevalid    => open                                                                        --               (terminated)
		);

	cpu_to_sdram_pb_m0_translator : component sopc_system_tse_dma_to_sdram_ccb_m0_translator
		generic map (
			AV_ADDRESS_W                => 27,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 27,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 1,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => sdram_0_afi_clk_clk,                                                   --                       clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                    --                     reset.reset
			uav_address              => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_to_sdram_pb_m0_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_to_sdram_pb_m0_waitrequest,                                        --                          .waitrequest
			av_burstcount            => cpu_to_sdram_pb_m0_burstcount,                                         --                          .burstcount
			av_byteenable            => cpu_to_sdram_pb_m0_byteenable,                                         --                          .byteenable
			av_read                  => cpu_to_sdram_pb_m0_read,                                               --                          .read
			av_readdata              => cpu_to_sdram_pb_m0_readdata,                                           --                          .readdata
			av_readdatavalid         => cpu_to_sdram_pb_m0_readdatavalid,                                      --                          .readdatavalid
			av_write                 => cpu_to_sdram_pb_m0_write,                                              --                          .write
			av_writedata             => cpu_to_sdram_pb_m0_writedata,                                          --                          .writedata
			av_debugaccess           => cpu_to_sdram_pb_m0_debugaccess,                                        --                          .debugaccess
			av_beginbursttransfer    => '0',                                                                   --               (terminated)
			av_begintransfer         => '0',                                                                   --               (terminated)
			av_chipselect            => '0',                                                                   --               (terminated)
			av_lock                  => '0',                                                                   --               (terminated)
			uav_clken                => open,                                                                  --               (terminated)
			av_clken                 => '1',                                                                   --               (terminated)
			uav_response             => "00",                                                                  --               (terminated)
			av_response              => open,                                                                  --               (terminated)
			uav_writeresponserequest => open,                                                                  --               (terminated)
			uav_writeresponsevalid   => '0',                                                                   --               (terminated)
			av_writeresponserequest  => '0',                                                                   --               (terminated)
			av_writeresponsevalid    => open                                                                   --               (terminated)
		);

	sdram_0_avl_translator : component sopc_system_sdram_0_avl_translator
		generic map (
			AV_ADDRESS_W                   => 24,
			AV_DATA_W                      => 64,
			UAV_DATA_W                     => 64,
			AV_BURSTCOUNT_W                => 3,
			AV_BYTEENABLE_W                => 8,
			UAV_BYTEENABLE_W               => 8,
			UAV_ADDRESS_W                  => 27,
			UAV_BURSTCOUNT_W               => 6,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 8,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_clk_clk,                                                    --                      clk.clk
			reset                    => rst_controller_004_reset_out_reset,                                     --                    reset.reset
			uav_address              => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sdram_0_avl_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sdram_0_avl_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => sdram_0_avl_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => sdram_0_avl_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sdram_0_avl_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_beginbursttransfer    => sdram_0_avl_translator_avalon_anti_slave_0_beginbursttransfer,          --                         .beginbursttransfer
			av_burstcount            => sdram_0_avl_translator_avalon_anti_slave_0_burstcount,                  --                         .burstcount
			av_byteenable            => sdram_0_avl_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => sdram_0_avl_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => sdram_0_avl_translator_avalon_anti_slave_0_inv,                         --                         .waitrequest
			av_begintransfer         => open,                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                   --              (terminated)
			av_lock                  => open,                                                                   --              (terminated)
			av_chipselect            => open,                                                                   --              (terminated)
			av_clken                 => open,                                                                   --              (terminated)
			uav_clken                => '0',                                                                    --              (terminated)
			av_debugaccess           => open,                                                                   --              (terminated)
			av_outputenable          => open,                                                                   --              (terminated)
			uav_response             => open,                                                                   --              (terminated)
			av_response              => "00",                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                     --              (terminated)
		);

	linux_cpu_tightly_coupled_data_master_0_translator : component sopc_system_linux_cpu_tightly_coupled_data_master_0_translator
		generic map (
			AV_ADDRESS_W                => 29,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 29,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => sdram_0_afi_clk_clk,                                                                        --                       clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                         --                     reset.reset
			uav_address              => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			uav_clken                => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_clken,         --                          .clken
			av_address               => linux_cpu_tightly_coupled_data_master_0_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => linux_cpu_tightly_coupled_data_master_0_waitrequest,                                        --                          .waitrequest
			av_byteenable            => linux_cpu_tightly_coupled_data_master_0_byteenable,                                         --                          .byteenable
			av_read                  => linux_cpu_tightly_coupled_data_master_0_read,                                               --                          .read
			av_readdata              => linux_cpu_tightly_coupled_data_master_0_readdata,                                           --                          .readdata
			av_readdatavalid         => linux_cpu_tightly_coupled_data_master_0_readdatavalid,                                      --                          .readdatavalid
			av_write                 => linux_cpu_tightly_coupled_data_master_0_write,                                              --                          .write
			av_writedata             => linux_cpu_tightly_coupled_data_master_0_writedata,                                          --                          .writedata
			av_clken                 => linux_cpu_tightly_coupled_data_master_0_clken,                                              --                          .clken
			av_burstcount            => "1",                                                                                        --               (terminated)
			av_beginbursttransfer    => '0',                                                                                        --               (terminated)
			av_begintransfer         => '0',                                                                                        --               (terminated)
			av_chipselect            => '0',                                                                                        --               (terminated)
			av_lock                  => '0',                                                                                        --               (terminated)
			av_debugaccess           => '0',                                                                                        --               (terminated)
			uav_response             => "00",                                                                                       --               (terminated)
			av_response              => open,                                                                                       --               (terminated)
			uav_writeresponserequest => open,                                                                                       --               (terminated)
			uav_writeresponsevalid   => '0',                                                                                        --               (terminated)
			av_writeresponserequest  => '0',                                                                                        --               (terminated)
			av_writeresponsevalid    => open                                                                                        --               (terminated)
		);

	tlb_miss_ram_1k_s1_translator : component sopc_system_tlb_miss_ram_1k_s1_translator
		generic map (
			AV_ADDRESS_W                   => 8,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 29,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 1,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_clk_clk,                                                                        --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                         --                    reset.reset
			uav_address              => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_burstcount,    --                         .burstcount
			uav_read                 => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_read,          --                         .read
			uav_write                => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_write,         --                         .write
			uav_waitrequest          => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_byteenable,    --                         .byteenable
			uav_readdata             => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_readdata,      --                         .readdata
			uav_writedata            => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_writedata,     --                         .writedata
			uav_lock                 => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_lock,          --                         .lock
			uav_debugaccess          => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_debugaccess,   --                         .debugaccess
			uav_clken                => linux_cpu_tightly_coupled_data_master_0_translator_avalon_universal_master_0_clken,         --                         .clken
			av_address               => tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_address,                                  --      avalon_anti_slave_0.address
			av_write                 => tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_write,                                    --                         .write
			av_readdata              => tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_readdata,                                 --                         .readdata
			av_writedata             => tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_writedata,                                --                         .writedata
			av_byteenable            => tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_byteenable,                               --                         .byteenable
			av_chipselect            => tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_chipselect,                               --                         .chipselect
			av_clken                 => tlb_miss_ram_1k_s1_translator_avalon_anti_slave_0_clken,                                    --                         .clken
			av_read                  => open,                                                                                       --              (terminated)
			av_begintransfer         => open,                                                                                       --              (terminated)
			av_beginbursttransfer    => open,                                                                                       --              (terminated)
			av_burstcount            => open,                                                                                       --              (terminated)
			av_readdatavalid         => '0',                                                                                        --              (terminated)
			av_waitrequest           => '0',                                                                                        --              (terminated)
			av_writebyteenable       => open,                                                                                       --              (terminated)
			av_lock                  => open,                                                                                       --              (terminated)
			av_debugaccess           => open,                                                                                       --              (terminated)
			av_outputenable          => open,                                                                                       --              (terminated)
			uav_response             => open,                                                                                       --              (terminated)
			av_response              => "00",                                                                                       --              (terminated)
			uav_writeresponserequest => '0',                                                                                        --              (terminated)
			uav_writeresponsevalid   => open,                                                                                       --              (terminated)
			av_writeresponserequest  => open,                                                                                       --              (terminated)
			av_writeresponsevalid    => '0'                                                                                         --              (terminated)
		);

	linux_cpu_tightly_coupled_instruction_master_0_translator : component sopc_system_linux_cpu_tightly_coupled_instruction_master_0_translator
		generic map (
			AV_ADDRESS_W                => 29,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 29,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => sdram_0_afi_clk_clk,                                                                               --                       clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                                --                     reset.reset
			uav_address              => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			uav_clken                => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_clken,         --                          .clken
			av_address               => linux_cpu_tightly_coupled_instruction_master_0_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => linux_cpu_tightly_coupled_instruction_master_0_waitrequest,                                        --                          .waitrequest
			av_read                  => linux_cpu_tightly_coupled_instruction_master_0_read,                                               --                          .read
			av_readdata              => linux_cpu_tightly_coupled_instruction_master_0_readdata,                                           --                          .readdata
			av_readdatavalid         => linux_cpu_tightly_coupled_instruction_master_0_readdatavalid,                                      --                          .readdatavalid
			av_clken                 => linux_cpu_tightly_coupled_instruction_master_0_clken,                                              --                          .clken
			av_burstcount            => "1",                                                                                               --               (terminated)
			av_byteenable            => "1111",                                                                                            --               (terminated)
			av_beginbursttransfer    => '0',                                                                                               --               (terminated)
			av_begintransfer         => '0',                                                                                               --               (terminated)
			av_chipselect            => '0',                                                                                               --               (terminated)
			av_write                 => '0',                                                                                               --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                                                --               (terminated)
			av_lock                  => '0',                                                                                               --               (terminated)
			av_debugaccess           => '0',                                                                                               --               (terminated)
			uav_response             => "00",                                                                                              --               (terminated)
			av_response              => open,                                                                                              --               (terminated)
			uav_writeresponserequest => open,                                                                                              --               (terminated)
			uav_writeresponsevalid   => '0',                                                                                               --               (terminated)
			av_writeresponserequest  => '0',                                                                                               --               (terminated)
			av_writeresponsevalid    => open                                                                                               --               (terminated)
		);

	tlb_miss_ram_1k_s2_translator : component sopc_system_tlb_miss_ram_1k_s1_translator
		generic map (
			AV_ADDRESS_W                   => 8,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 29,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 1,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => sdram_0_afi_clk_clk,                                                                               --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                                --                    reset.reset
			uav_address              => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_burstcount,    --                         .burstcount
			uav_read                 => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_read,          --                         .read
			uav_write                => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_write,         --                         .write
			uav_waitrequest          => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_byteenable,    --                         .byteenable
			uav_readdata             => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_readdata,      --                         .readdata
			uav_writedata            => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_writedata,     --                         .writedata
			uav_lock                 => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_lock,          --                         .lock
			uav_debugaccess          => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_debugaccess,   --                         .debugaccess
			uav_clken                => linux_cpu_tightly_coupled_instruction_master_0_translator_avalon_universal_master_0_clken,         --                         .clken
			av_address               => tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_address,                                         --      avalon_anti_slave_0.address
			av_write                 => tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_write,                                           --                         .write
			av_readdata              => tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_readdata,                                        --                         .readdata
			av_writedata             => tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_writedata,                                       --                         .writedata
			av_byteenable            => tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_byteenable,                                      --                         .byteenable
			av_chipselect            => tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_chipselect,                                      --                         .chipselect
			av_clken                 => tlb_miss_ram_1k_s2_translator_avalon_anti_slave_0_clken,                                           --                         .clken
			av_read                  => open,                                                                                              --              (terminated)
			av_begintransfer         => open,                                                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                                                              --              (terminated)
			av_burstcount            => open,                                                                                              --              (terminated)
			av_readdatavalid         => '0',                                                                                               --              (terminated)
			av_waitrequest           => '0',                                                                                               --              (terminated)
			av_writebyteenable       => open,                                                                                              --              (terminated)
			av_lock                  => open,                                                                                              --              (terminated)
			av_debugaccess           => open,                                                                                              --              (terminated)
			av_outputenable          => open,                                                                                              --              (terminated)
			uav_response             => open,                                                                                              --              (terminated)
			av_response              => "00",                                                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                                                              --              (terminated)
			av_writeresponserequest  => open,                                                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                                                --              (terminated)
		);

	linux_cpu_data_master_translator_avalon_universal_master_0_agent : component sopc_system_linux_cpu_data_master_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_BEGIN_BURST           => 84,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 74,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			PKT_BURST_TYPE_H          => 81,
			PKT_BURST_TYPE_L          => 80,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_ADDR_H                => 64,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 65,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			PKT_TRANS_READ            => 68,
			PKT_TRANS_LOCK            => 69,
			PKT_TRANS_EXCLUSIVE       => 70,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 88,
			PKT_THREAD_ID_H           => 90,
			PKT_THREAD_ID_L           => 90,
			PKT_CACHE_H               => 97,
			PKT_CACHE_L               => 94,
			PKT_DATA_SIDEBAND_H       => 83,
			PKT_DATA_SIDEBAND_L       => 83,
			PKT_QOS_H                 => 85,
			PKT_QOS_L                 => 85,
			PKT_ADDR_SIDEBAND_H       => 82,
			PKT_ADDR_SIDEBAND_L       => 82,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			ST_DATA_W                 => 100,
			ST_CHANNEL_W              => 4,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_clk_clk,                                                               --       clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                -- clk_reset.reset
			av_address              => linux_cpu_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => linux_cpu_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => linux_cpu_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => linux_cpu_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => linux_cpu_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => linux_cpu_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => linux_cpu_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => linux_cpu_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => linux_cpu_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => linux_cpu_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => linux_cpu_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => linux_cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => linux_cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => linux_cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => linux_cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => linux_cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => limiter_rsp_src_valid,                                                             --        rp.valid
			rp_data                 => limiter_rsp_src_data,                                                              --          .data
			rp_channel              => limiter_rsp_src_channel,                                                           --          .channel
			rp_startofpacket        => limiter_rsp_src_startofpacket,                                                     --          .startofpacket
			rp_endofpacket          => limiter_rsp_src_endofpacket,                                                       --          .endofpacket
			rp_ready                => limiter_rsp_src_ready,                                                             --          .ready
			av_response             => open,                                                                              -- (terminated)
			av_writeresponserequest => '0',                                                                               -- (terminated)
			av_writeresponsevalid   => open                                                                               -- (terminated)
		);

	linux_cpu_instruction_master_translator_avalon_universal_master_0_agent : component sopc_system_linux_cpu_data_master_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_BEGIN_BURST           => 84,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 74,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			PKT_BURST_TYPE_H          => 81,
			PKT_BURST_TYPE_L          => 80,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_ADDR_H                => 64,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 65,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			PKT_TRANS_READ            => 68,
			PKT_TRANS_LOCK            => 69,
			PKT_TRANS_EXCLUSIVE       => 70,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 88,
			PKT_THREAD_ID_H           => 90,
			PKT_THREAD_ID_L           => 90,
			PKT_CACHE_H               => 97,
			PKT_CACHE_L               => 94,
			PKT_DATA_SIDEBAND_H       => 83,
			PKT_DATA_SIDEBAND_L       => 83,
			PKT_QOS_H                 => 85,
			PKT_QOS_L                 => 85,
			PKT_ADDR_SIDEBAND_H       => 82,
			PKT_ADDR_SIDEBAND_L       => 82,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			ST_DATA_W                 => 100,
			ST_CHANNEL_W              => 4,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 3,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_clk_clk,                                                                      --       clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                       -- clk_reset.reset
			av_address              => linux_cpu_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => linux_cpu_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => linux_cpu_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => linux_cpu_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => linux_cpu_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => linux_cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => linux_cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => linux_cpu_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => linux_cpu_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => linux_cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => linux_cpu_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => linux_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => linux_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => linux_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => linux_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => linux_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => limiter_001_rsp_src_valid,                                                                --        rp.valid
			rp_data                 => limiter_001_rsp_src_data,                                                                 --          .data
			rp_channel              => limiter_001_rsp_src_channel,                                                              --          .channel
			rp_startofpacket        => limiter_001_rsp_src_startofpacket,                                                        --          .startofpacket
			rp_endofpacket          => limiter_001_rsp_src_endofpacket,                                                          --          .endofpacket
			rp_ready                => limiter_001_rsp_src_ready,                                                                --          .ready
			av_response             => open,                                                                                     -- (terminated)
			av_writeresponserequest => '0',                                                                                      -- (terminated)
			av_writeresponsevalid   => open                                                                                      -- (terminated)
		);

	linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent : component sopc_system_linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 84,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 64,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 65,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			PKT_TRANS_READ            => 68,
			PKT_TRANS_LOCK            => 69,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 74,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			ST_CHANNEL_W              => 4,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_clk_clk,                                                                              --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                               --       clk_reset.reset
			m0_address              => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_src_ready,                                                                           --              cp.ready
			cp_valid                => cmd_xbar_mux_src_valid,                                                                           --                .valid
			cp_data                 => cmd_xbar_mux_src_data,                                                                            --                .data
			cp_startofpacket        => cmd_xbar_mux_src_startofpacket,                                                                   --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_src_endofpacket,                                                                     --                .endofpacket
			cp_channel              => cmd_xbar_mux_src_channel,                                                                         --                .channel
			rf_sink_ready           => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                               --     (terminated)
		);

	linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_clk_clk,                                                                              --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                               -- clk_reset.reset
			in_data           => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                             -- (terminated)
			csr_read          => '0',                                                                                              -- (terminated)
			csr_write         => '0',                                                                                              -- (terminated)
			csr_readdata      => open,                                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                               -- (terminated)
			almost_full_data  => open,                                                                                             -- (terminated)
			almost_empty_data => open,                                                                                             -- (terminated)
			in_empty          => '0',                                                                                              -- (terminated)
			out_empty         => open,                                                                                             -- (terminated)
			in_error          => '0',                                                                                              -- (terminated)
			out_error         => open,                                                                                             -- (terminated)
			in_channel        => '0',                                                                                              -- (terminated)
			out_channel       => open                                                                                              -- (terminated)
		);

	cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent : component sopc_system_linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 84,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 64,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 65,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			PKT_TRANS_READ            => 68,
			PKT_TRANS_LOCK            => 69,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 74,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			ST_CHANNEL_W              => 4,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_clk_clk,                                                                      --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                       --       clk_reset.reset
			m0_address              => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_001_src_ready,                                                               --              cp.ready
			cp_valid                => cmd_xbar_mux_001_src_valid,                                                               --                .valid
			cp_data                 => cmd_xbar_mux_001_src_data,                                                                --                .data
			cp_startofpacket        => cmd_xbar_mux_001_src_startofpacket,                                                       --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_001_src_endofpacket,                                                         --                .endofpacket
			cp_channel              => cmd_xbar_mux_001_src_channel,                                                             --                .channel
			rf_sink_ready           => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                     --     (terminated)
			m0_writeresponserequest => open,                                                                                     --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                       --     (terminated)
		);

	cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 9,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_clk_clk,                                                                      --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                       -- clk_reset.reset
			in_data           => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                     -- (terminated)
			csr_read          => '0',                                                                                      -- (terminated)
			csr_write         => '0',                                                                                      -- (terminated)
			csr_readdata      => open,                                                                                     -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                       -- (terminated)
			almost_full_data  => open,                                                                                     -- (terminated)
			almost_empty_data => open,                                                                                     -- (terminated)
			in_empty          => '0',                                                                                      -- (terminated)
			out_empty         => open,                                                                                     -- (terminated)
			in_error          => '0',                                                                                      -- (terminated)
			out_error         => open,                                                                                     -- (terminated)
			in_channel        => '0',                                                                                      -- (terminated)
			out_channel       => open                                                                                      -- (terminated)
		);

	cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent : component sopc_system_linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 84,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 64,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 65,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			PKT_TRANS_READ            => 68,
			PKT_TRANS_LOCK            => 69,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 74,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			ST_CHANNEL_W              => 4,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_clk_clk,                                                                            --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                             --       clk_reset.reset
			m0_address              => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_src2_ready,                                                                      --              cp.ready
			cp_valid                => cmd_xbar_demux_src2_valid,                                                                      --                .valid
			cp_data                 => cmd_xbar_demux_src2_data,                                                                       --                .data
			cp_startofpacket        => cmd_xbar_demux_src2_startofpacket,                                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_src2_endofpacket,                                                                --                .endofpacket
			cp_channel              => cmd_xbar_demux_src2_channel,                                                                    --                .channel
			rf_sink_ready           => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                             --     (terminated)
		);

	cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 9,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_clk_clk,                                                                            --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                             -- clk_reset.reset
			in_data           => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                           -- (terminated)
			csr_read          => '0',                                                                                            -- (terminated)
			csr_write         => '0',                                                                                            -- (terminated)
			csr_readdata      => open,                                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                             -- (terminated)
			almost_full_data  => open,                                                                                           -- (terminated)
			almost_empty_data => open,                                                                                           -- (terminated)
			in_empty          => '0',                                                                                            -- (terminated)
			out_empty         => open,                                                                                           -- (terminated)
			in_error          => '0',                                                                                            -- (terminated)
			out_error         => open,                                                                                           -- (terminated)
			in_channel        => '0',                                                                                            -- (terminated)
			out_channel       => open                                                                                            -- (terminated)
		);

	cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent : component sopc_system_linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 84,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 64,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 65,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			PKT_TRANS_READ            => 68,
			PKT_TRANS_LOCK            => 69,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 86,
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 76,
			PKT_BURSTWRAP_L           => 74,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_PROTECTION_H          => 93,
			PKT_PROTECTION_L          => 91,
			PKT_RESPONSE_STATUS_H     => 99,
			PKT_RESPONSE_STATUS_L     => 98,
			PKT_BURST_SIZE_H          => 79,
			PKT_BURST_SIZE_L          => 77,
			ST_CHANNEL_W              => 4,
			ST_DATA_W                 => 100,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_clk_clk,                                                                     --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                      --       clk_reset.reset
			m0_address              => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_003_src_ready,                                                              --              cp.ready
			cp_valid                => cmd_xbar_mux_003_src_valid,                                                              --                .valid
			cp_data                 => cmd_xbar_mux_003_src_data,                                                               --                .data
			cp_startofpacket        => cmd_xbar_mux_003_src_startofpacket,                                                      --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_003_src_endofpacket,                                                        --                .endofpacket
			cp_channel              => cmd_xbar_mux_003_src_channel,                                                            --                .channel
			rf_sink_ready           => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                    --     (terminated)
			m0_writeresponserequest => open,                                                                                    --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                      --     (terminated)
		);

	cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 101,
			FIFO_DEPTH          => 5,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_clk_clk,                                                                     --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                      -- clk_reset.reset
			in_data           => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                    -- (terminated)
			csr_read          => '0',                                                                                     -- (terminated)
			csr_write         => '0',                                                                                     -- (terminated)
			csr_readdata      => open,                                                                                    -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                      -- (terminated)
			almost_full_data  => open,                                                                                    -- (terminated)
			almost_empty_data => open,                                                                                    -- (terminated)
			in_empty          => '0',                                                                                     -- (terminated)
			out_empty         => open,                                                                                    -- (terminated)
			in_error          => '0',                                                                                     -- (terminated)
			out_error         => open,                                                                                    -- (terminated)
			in_channel        => '0',                                                                                     -- (terminated)
			out_channel       => open                                                                                     -- (terminated)
		);

	sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent : component sopc_system_sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 94,
			PKT_PROTECTION_L          => 92,
			PKT_BEGIN_BURST           => 85,
			PKT_BURSTWRAP_H           => 77,
			PKT_BURSTWRAP_L           => 77,
			PKT_BURST_SIZE_H          => 80,
			PKT_BURST_SIZE_L          => 78,
			PKT_BURST_TYPE_H          => 82,
			PKT_BURST_TYPE_L          => 81,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 88,
			PKT_SRC_ID_L              => 87,
			PKT_DEST_ID_H             => 90,
			PKT_DEST_ID_L             => 89,
			PKT_THREAD_ID_H           => 91,
			PKT_THREAD_ID_L           => 91,
			PKT_CACHE_H               => 98,
			PKT_CACHE_L               => 95,
			PKT_DATA_SIDEBAND_H       => 84,
			PKT_DATA_SIDEBAND_L       => 84,
			PKT_QOS_H                 => 86,
			PKT_QOS_L                 => 86,
			PKT_ADDR_SIDEBAND_H       => 83,
			PKT_ADDR_SIDEBAND_L       => 83,
			PKT_RESPONSE_STATUS_H     => 100,
			PKT_RESPONSE_STATUS_L     => 99,
			ST_DATA_W                 => 101,
			ST_CHANNEL_W              => 4,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 3,
			BURSTWRAP_VALUE           => 1,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                              --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			av_address              => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_demux_004_src0_valid,                                                         --        rp.valid
			rp_data                 => rsp_xbar_demux_004_src0_data,                                                          --          .data
			rp_channel              => rsp_xbar_demux_004_src0_channel,                                                       --          .channel
			rp_startofpacket        => rsp_xbar_demux_004_src0_startofpacket,                                                 --          .startofpacket
			rp_endofpacket          => rsp_xbar_demux_004_src0_endofpacket,                                                   --          .endofpacket
			rp_ready                => rsp_xbar_demux_004_src0_ready,                                                         --          .ready
			av_response             => open,                                                                                  -- (terminated)
			av_writeresponserequest => '0',                                                                                   -- (terminated)
			av_writeresponsevalid   => open                                                                                   -- (terminated)
		);

	sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent : component sopc_system_sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 94,
			PKT_PROTECTION_L          => 92,
			PKT_BEGIN_BURST           => 85,
			PKT_BURSTWRAP_H           => 77,
			PKT_BURSTWRAP_L           => 77,
			PKT_BURST_SIZE_H          => 80,
			PKT_BURST_SIZE_L          => 78,
			PKT_BURST_TYPE_H          => 82,
			PKT_BURST_TYPE_L          => 81,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 88,
			PKT_SRC_ID_L              => 87,
			PKT_DEST_ID_H             => 90,
			PKT_DEST_ID_L             => 89,
			PKT_THREAD_ID_H           => 91,
			PKT_THREAD_ID_L           => 91,
			PKT_CACHE_H               => 98,
			PKT_CACHE_L               => 95,
			PKT_DATA_SIDEBAND_H       => 84,
			PKT_DATA_SIDEBAND_L       => 84,
			PKT_QOS_H                 => 86,
			PKT_QOS_L                 => 86,
			PKT_ADDR_SIDEBAND_H       => 83,
			PKT_ADDR_SIDEBAND_L       => 83,
			PKT_RESPONSE_STATUS_H     => 100,
			PKT_RESPONSE_STATUS_L     => 99,
			ST_DATA_W                 => 101,
			ST_CHANNEL_W              => 4,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 1,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                              --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			av_address              => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_demux_004_src1_valid,                                                         --        rp.valid
			rp_data                 => rsp_xbar_demux_004_src1_data,                                                          --          .data
			rp_channel              => rsp_xbar_demux_004_src1_channel,                                                       --          .channel
			rp_startofpacket        => rsp_xbar_demux_004_src1_startofpacket,                                                 --          .startofpacket
			rp_endofpacket          => rsp_xbar_demux_004_src1_endofpacket,                                                   --          .endofpacket
			rp_ready                => rsp_xbar_demux_004_src1_ready,                                                         --          .ready
			av_response             => open,                                                                                  -- (terminated)
			av_writeresponserequest => '0',                                                                                   -- (terminated)
			av_writeresponsevalid   => open                                                                                   -- (terminated)
		);

	sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent : component sopc_system_sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 94,
			PKT_PROTECTION_L          => 92,
			PKT_BEGIN_BURST           => 85,
			PKT_BURSTWRAP_H           => 77,
			PKT_BURSTWRAP_L           => 77,
			PKT_BURST_SIZE_H          => 80,
			PKT_BURST_SIZE_L          => 78,
			PKT_BURST_TYPE_H          => 82,
			PKT_BURST_TYPE_L          => 81,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 88,
			PKT_SRC_ID_L              => 87,
			PKT_DEST_ID_H             => 90,
			PKT_DEST_ID_L             => 89,
			PKT_THREAD_ID_H           => 91,
			PKT_THREAD_ID_L           => 91,
			PKT_CACHE_H               => 98,
			PKT_CACHE_L               => 95,
			PKT_DATA_SIDEBAND_H       => 84,
			PKT_DATA_SIDEBAND_L       => 84,
			PKT_QOS_H                 => 86,
			PKT_QOS_L                 => 86,
			PKT_ADDR_SIDEBAND_H       => 83,
			PKT_ADDR_SIDEBAND_L       => 83,
			PKT_RESPONSE_STATUS_H     => 100,
			PKT_RESPONSE_STATUS_L     => 99,
			ST_DATA_W                 => 101,
			ST_CHANNEL_W              => 4,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 1,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                             --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			av_address              => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_demux_004_src2_valid,                                                        --        rp.valid
			rp_data                 => rsp_xbar_demux_004_src2_data,                                                         --          .data
			rp_channel              => rsp_xbar_demux_004_src2_channel,                                                      --          .channel
			rp_startofpacket        => rsp_xbar_demux_004_src2_startofpacket,                                                --          .startofpacket
			rp_endofpacket          => rsp_xbar_demux_004_src2_endofpacket,                                                  --          .endofpacket
			rp_ready                => rsp_xbar_demux_004_src2_ready,                                                        --          .ready
			av_response             => open,                                                                                 -- (terminated)
			av_writeresponserequest => '0',                                                                                  -- (terminated)
			av_writeresponsevalid   => open                                                                                  -- (terminated)
		);

	sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent : component sopc_system_sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 94,
			PKT_PROTECTION_L          => 92,
			PKT_BEGIN_BURST           => 85,
			PKT_BURSTWRAP_H           => 77,
			PKT_BURSTWRAP_L           => 77,
			PKT_BURST_SIZE_H          => 80,
			PKT_BURST_SIZE_L          => 78,
			PKT_BURST_TYPE_H          => 82,
			PKT_BURST_TYPE_L          => 81,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 88,
			PKT_SRC_ID_L              => 87,
			PKT_DEST_ID_H             => 90,
			PKT_DEST_ID_L             => 89,
			PKT_THREAD_ID_H           => 91,
			PKT_THREAD_ID_L           => 91,
			PKT_CACHE_H               => 98,
			PKT_CACHE_L               => 95,
			PKT_DATA_SIDEBAND_H       => 84,
			PKT_DATA_SIDEBAND_L       => 84,
			PKT_QOS_H                 => 86,
			PKT_QOS_L                 => 86,
			PKT_ADDR_SIDEBAND_H       => 83,
			PKT_ADDR_SIDEBAND_L       => 83,
			PKT_RESPONSE_STATUS_H     => 100,
			PKT_RESPONSE_STATUS_L     => 99,
			ST_DATA_W                 => 101,
			ST_CHANNEL_W              => 4,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 2,
			BURSTWRAP_VALUE           => 1,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                             --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			av_address              => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_demux_004_src3_valid,                                                        --        rp.valid
			rp_data                 => rsp_xbar_demux_004_src3_data,                                                         --          .data
			rp_channel              => rsp_xbar_demux_004_src3_channel,                                                      --          .channel
			rp_startofpacket        => rsp_xbar_demux_004_src3_startofpacket,                                                --          .startofpacket
			rp_endofpacket          => rsp_xbar_demux_004_src3_endofpacket,                                                  --          .endofpacket
			rp_ready                => rsp_xbar_demux_004_src3_ready,                                                        --          .ready
			av_response             => open,                                                                                 -- (terminated)
			av_writeresponserequest => '0',                                                                                  -- (terminated)
			av_writeresponsevalid   => open                                                                                  -- (terminated)
		);

	dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent : component sopc_system_dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 85,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 88,
			PKT_SRC_ID_L              => 87,
			PKT_DEST_ID_H             => 90,
			PKT_DEST_ID_L             => 89,
			PKT_BURSTWRAP_H           => 77,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 94,
			PKT_PROTECTION_L          => 92,
			PKT_RESPONSE_STATUS_H     => 100,
			PKT_RESPONSE_STATUS_L     => 99,
			PKT_BURST_SIZE_H          => 80,
			PKT_BURST_SIZE_L          => 78,
			ST_CHANNEL_W              => 4,
			ST_DATA_W                 => 101,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                                      --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                --       clk_reset.reset
			m0_address              => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_004_src_ready,                                                                    --              cp.ready
			cp_valid                => cmd_xbar_mux_004_src_valid,                                                                    --                .valid
			cp_data                 => cmd_xbar_mux_004_src_data,                                                                     --                .data
			cp_startofpacket        => cmd_xbar_mux_004_src_startofpacket,                                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_004_src_endofpacket,                                                              --                .endofpacket
			cp_channel              => cmd_xbar_mux_004_src_channel,                                                                  --                .channel
			rf_sink_ready           => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                          --     (terminated)
			m0_writeresponserequest => open,                                                                                          --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                            --     (terminated)
		);

	dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 102,
			FIFO_DEPTH          => 5,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_half_clk_clk,                                                                      --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                -- clk_reset.reset
			in_data           => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                          -- (terminated)
			csr_read          => '0',                                                                                           -- (terminated)
			csr_write         => '0',                                                                                           -- (terminated)
			csr_readdata      => open,                                                                                          -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                            -- (terminated)
			almost_full_data  => open,                                                                                          -- (terminated)
			almost_empty_data => open,                                                                                          -- (terminated)
			in_empty          => '0',                                                                                           -- (terminated)
			out_empty         => open,                                                                                          -- (terminated)
			in_error          => '0',                                                                                           -- (terminated)
			out_error         => open,                                                                                          -- (terminated)
			in_channel        => '0',                                                                                           -- (terminated)
			out_channel       => open                                                                                           -- (terminated)
		);

	dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent : component sopc_system_dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 87,
			PKT_PROTECTION_L          => 85,
			PKT_BEGIN_BURST           => 76,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 68,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			PKT_BURST_TYPE_H          => 73,
			PKT_BURST_TYPE_L          => 72,
			PKT_BYTE_CNT_H            => 67,
			PKT_BYTE_CNT_L            => 65,
			PKT_ADDR_H                => 58,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 59,
			PKT_TRANS_POSTED          => 60,
			PKT_TRANS_WRITE           => 61,
			PKT_TRANS_READ            => 62,
			PKT_TRANS_LOCK            => 63,
			PKT_TRANS_EXCLUSIVE       => 64,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 83,
			PKT_DEST_ID_L             => 81,
			PKT_THREAD_ID_H           => 84,
			PKT_THREAD_ID_L           => 84,
			PKT_CACHE_H               => 91,
			PKT_CACHE_L               => 88,
			PKT_DATA_SIDEBAND_H       => 75,
			PKT_DATA_SIDEBAND_L       => 75,
			PKT_QOS_H                 => 77,
			PKT_QOS_L                 => 77,
			PKT_ADDR_SIDEBAND_H       => 74,
			PKT_ADDR_SIDEBAND_L       => 74,
			PKT_RESPONSE_STATUS_H     => 93,
			PKT_RESPONSE_STATUS_L     => 92,
			ST_DATA_W                 => 94,
			ST_CHANNEL_W              => 8,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 1,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                             --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			av_address              => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_demux_005_src0_valid,                                                        --        rp.valid
			rp_data                 => rsp_xbar_demux_005_src0_data,                                                         --          .data
			rp_channel              => rsp_xbar_demux_005_src0_channel,                                                      --          .channel
			rp_startofpacket        => rsp_xbar_demux_005_src0_startofpacket,                                                --          .startofpacket
			rp_endofpacket          => rsp_xbar_demux_005_src0_endofpacket,                                                  --          .endofpacket
			rp_ready                => rsp_xbar_demux_005_src0_ready,                                                        --          .ready
			av_response             => open,                                                                                 -- (terminated)
			av_writeresponserequest => '0',                                                                                  -- (terminated)
			av_writeresponsevalid   => open                                                                                  -- (terminated)
		);

	cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent : component sopc_system_dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 87,
			PKT_PROTECTION_L          => 85,
			PKT_BEGIN_BURST           => 76,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 68,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			PKT_BURST_TYPE_H          => 73,
			PKT_BURST_TYPE_L          => 72,
			PKT_BYTE_CNT_H            => 67,
			PKT_BYTE_CNT_L            => 65,
			PKT_ADDR_H                => 58,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 59,
			PKT_TRANS_POSTED          => 60,
			PKT_TRANS_WRITE           => 61,
			PKT_TRANS_READ            => 62,
			PKT_TRANS_LOCK            => 63,
			PKT_TRANS_EXCLUSIVE       => 64,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 83,
			PKT_DEST_ID_L             => 81,
			PKT_THREAD_ID_H           => 84,
			PKT_THREAD_ID_L           => 84,
			PKT_CACHE_H               => 91,
			PKT_CACHE_L               => 88,
			PKT_DATA_SIDEBAND_H       => 75,
			PKT_DATA_SIDEBAND_L       => 75,
			PKT_QOS_H                 => 77,
			PKT_QOS_L                 => 77,
			PKT_ADDR_SIDEBAND_H       => 74,
			PKT_ADDR_SIDEBAND_L       => 74,
			PKT_RESPONSE_STATUS_H     => 93,
			PKT_RESPONSE_STATUS_L     => 92,
			ST_DATA_W                 => 94,
			ST_CHANNEL_W              => 8,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 1,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                              --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			av_address              => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => limiter_002_rsp_src_valid,                                                             --        rp.valid
			rp_data                 => limiter_002_rsp_src_data,                                                              --          .data
			rp_channel              => limiter_002_rsp_src_channel,                                                           --          .channel
			rp_startofpacket        => limiter_002_rsp_src_startofpacket,                                                     --          .startofpacket
			rp_endofpacket          => limiter_002_rsp_src_endofpacket,                                                       --          .endofpacket
			rp_ready                => limiter_002_rsp_src_ready,                                                             --          .ready
			av_response             => open,                                                                                  -- (terminated)
			av_writeresponserequest => '0',                                                                                   -- (terminated)
			av_writeresponsevalid   => open                                                                                   -- (terminated)
		);

	descriptor_memory_s1_translator_avalon_universal_slave_0_agent : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 58,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 59,
			PKT_TRANS_POSTED          => 60,
			PKT_TRANS_WRITE           => 61,
			PKT_TRANS_READ            => 62,
			PKT_TRANS_LOCK            => 63,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 83,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 68,
			PKT_BYTE_CNT_H            => 67,
			PKT_BYTE_CNT_L            => 65,
			PKT_PROTECTION_H          => 87,
			PKT_PROTECTION_L          => 85,
			PKT_RESPONSE_STATUS_H     => 93,
			PKT_RESPONSE_STATUS_L     => 92,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 94,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                                  --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                            --       clk_reset.reset
			m0_address              => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_005_src_ready,                                                                --              cp.ready
			cp_valid                => cmd_xbar_mux_005_src_valid,                                                                --                .valid
			cp_data                 => cmd_xbar_mux_005_src_data,                                                                 --                .data
			cp_startofpacket        => cmd_xbar_mux_005_src_startofpacket,                                                        --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_005_src_endofpacket,                                                          --                .endofpacket
			cp_channel              => cmd_xbar_mux_005_src_channel,                                                              --                .channel
			rf_sink_ready           => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                      --     (terminated)
			m0_writeresponserequest => open,                                                                                      --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                        --     (terminated)
		);

	descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 95,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_half_clk_clk,                                                                  --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			in_data           => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                      -- (terminated)
			csr_read          => '0',                                                                                       -- (terminated)
			csr_write         => '0',                                                                                       -- (terminated)
			csr_readdata      => open,                                                                                      -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                        -- (terminated)
			almost_full_data  => open,                                                                                      -- (terminated)
			almost_empty_data => open,                                                                                      -- (terminated)
			in_empty          => '0',                                                                                       -- (terminated)
			out_empty         => open,                                                                                      -- (terminated)
			in_error          => '0',                                                                                       -- (terminated)
			out_error         => open,                                                                                      -- (terminated)
			in_channel        => '0',                                                                                       -- (terminated)
			out_channel       => open                                                                                       -- (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 58,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 59,
			PKT_TRANS_POSTED          => 60,
			PKT_TRANS_WRITE           => 61,
			PKT_TRANS_READ            => 62,
			PKT_TRANS_LOCK            => 63,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 83,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 68,
			PKT_BYTE_CNT_H            => 67,
			PKT_BYTE_CNT_L            => 65,
			PKT_PROTECTION_H          => 87,
			PKT_PROTECTION_L          => 85,
			PKT_RESPONSE_STATUS_H     => 93,
			PKT_RESPONSE_STATUS_L     => 92,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 94,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                   --       clk_reset.reset
			m0_address              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_007_src1_ready,                                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_007_src1_valid,                                                                    --                .valid
			cp_data                 => cmd_xbar_demux_007_src1_data,                                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_007_src1_startofpacket,                                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_007_src1_endofpacket,                                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_007_src1_channel,                                                                  --                .channel
			rf_sink_ready           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                               --     (terminated)
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 95,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_half_clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                   -- clk_reset.reset
			in_data           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                             -- (terminated)
			csr_read          => '0',                                                                                              -- (terminated)
			csr_write         => '0',                                                                                              -- (terminated)
			csr_readdata      => open,                                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                               -- (terminated)
			almost_full_data  => open,                                                                                             -- (terminated)
			almost_empty_data => open,                                                                                             -- (terminated)
			in_empty          => '0',                                                                                              -- (terminated)
			out_empty         => open,                                                                                             -- (terminated)
			in_error          => '0',                                                                                              -- (terminated)
			out_error         => open,                                                                                             -- (terminated)
			in_channel        => '0',                                                                                              -- (terminated)
			out_channel       => open                                                                                              -- (terminated)
		);

	tse_mac_control_port_translator_avalon_universal_slave_0_agent : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 58,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 59,
			PKT_TRANS_POSTED          => 60,
			PKT_TRANS_WRITE           => 61,
			PKT_TRANS_READ            => 62,
			PKT_TRANS_LOCK            => 63,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 83,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 68,
			PKT_BYTE_CNT_H            => 67,
			PKT_BYTE_CNT_L            => 65,
			PKT_PROTECTION_H          => 87,
			PKT_PROTECTION_L          => 85,
			PKT_RESPONSE_STATUS_H     => 93,
			PKT_RESPONSE_STATUS_L     => 92,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 94,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                                  --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                            --       clk_reset.reset
			m0_address              => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => tse_mac_control_port_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_007_src2_ready,                                                             --              cp.ready
			cp_valid                => cmd_xbar_demux_007_src2_valid,                                                             --                .valid
			cp_data                 => cmd_xbar_demux_007_src2_data,                                                              --                .data
			cp_startofpacket        => cmd_xbar_demux_007_src2_startofpacket,                                                     --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_007_src2_endofpacket,                                                       --                .endofpacket
			cp_channel              => cmd_xbar_demux_007_src2_channel,                                                           --                .channel
			rf_sink_ready           => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                      --     (terminated)
			m0_writeresponserequest => open,                                                                                      --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                        --     (terminated)
		);

	tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 95,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_half_clk_clk,                                                                  --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			in_data           => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                      -- (terminated)
			csr_read          => '0',                                                                                       -- (terminated)
			csr_write         => '0',                                                                                       -- (terminated)
			csr_readdata      => open,                                                                                      -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                        -- (terminated)
			almost_full_data  => open,                                                                                      -- (terminated)
			almost_empty_data => open,                                                                                      -- (terminated)
			in_empty          => '0',                                                                                       -- (terminated)
			out_empty         => open,                                                                                      -- (terminated)
			in_error          => '0',                                                                                       -- (terminated)
			out_error         => open,                                                                                      -- (terminated)
			in_channel        => '0',                                                                                       -- (terminated)
			out_channel       => open                                                                                       -- (terminated)
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 58,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 59,
			PKT_TRANS_POSTED          => 60,
			PKT_TRANS_WRITE           => 61,
			PKT_TRANS_READ            => 62,
			PKT_TRANS_LOCK            => 63,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 83,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 68,
			PKT_BYTE_CNT_H            => 67,
			PKT_BYTE_CNT_L            => 65,
			PKT_PROTECTION_H          => 87,
			PKT_PROTECTION_L          => 85,
			PKT_RESPONSE_STATUS_H     => 93,
			PKT_RESPONSE_STATUS_L     => 92,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 94,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                                 --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                           --       clk_reset.reset
			m0_address              => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_007_src3_ready,                                                            --              cp.ready
			cp_valid                => cmd_xbar_demux_007_src3_valid,                                                            --                .valid
			cp_data                 => cmd_xbar_demux_007_src3_data,                                                             --                .data
			cp_startofpacket        => cmd_xbar_demux_007_src3_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_007_src3_endofpacket,                                                      --                .endofpacket
			cp_channel              => cmd_xbar_demux_007_src3_channel,                                                          --                .channel
			rf_sink_ready           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                     --     (terminated)
			m0_writeresponserequest => open,                                                                                     --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                       --     (terminated)
		);

	sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 95,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_half_clk_clk,                                                                 --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                           -- clk_reset.reset
			in_data           => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                     -- (terminated)
			csr_read          => '0',                                                                                      -- (terminated)
			csr_write         => '0',                                                                                      -- (terminated)
			csr_readdata      => open,                                                                                     -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                       -- (terminated)
			almost_full_data  => open,                                                                                     -- (terminated)
			almost_empty_data => open,                                                                                     -- (terminated)
			in_empty          => '0',                                                                                      -- (terminated)
			out_empty         => open,                                                                                     -- (terminated)
			in_error          => '0',                                                                                      -- (terminated)
			out_error         => open,                                                                                     -- (terminated)
			in_channel        => '0',                                                                                      -- (terminated)
			out_channel       => open                                                                                      -- (terminated)
		);

	linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 58,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 59,
			PKT_TRANS_POSTED          => 60,
			PKT_TRANS_WRITE           => 61,
			PKT_TRANS_READ            => 62,
			PKT_TRANS_LOCK            => 63,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 83,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 68,
			PKT_BYTE_CNT_H            => 67,
			PKT_BYTE_CNT_L            => 65,
			PKT_PROTECTION_H          => 87,
			PKT_PROTECTION_L          => 85,
			PKT_RESPONSE_STATUS_H     => 93,
			PKT_RESPONSE_STATUS_L     => 92,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 94,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                                --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                          --       clk_reset.reset
			m0_address              => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_007_src4_ready,                                                           --              cp.ready
			cp_valid                => cmd_xbar_demux_007_src4_valid,                                                           --                .valid
			cp_data                 => cmd_xbar_demux_007_src4_data,                                                            --                .data
			cp_startofpacket        => cmd_xbar_demux_007_src4_startofpacket,                                                   --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_007_src4_endofpacket,                                                     --                .endofpacket
			cp_channel              => cmd_xbar_demux_007_src4_channel,                                                         --                .channel
			rf_sink_ready           => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                    --     (terminated)
			m0_writeresponserequest => open,                                                                                    --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                      --     (terminated)
		);

	linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 95,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_half_clk_clk,                                                                --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                          -- clk_reset.reset
			in_data           => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                    -- (terminated)
			csr_read          => '0',                                                                                     -- (terminated)
			csr_write         => '0',                                                                                     -- (terminated)
			csr_readdata      => open,                                                                                    -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                      -- (terminated)
			almost_full_data  => open,                                                                                    -- (terminated)
			almost_empty_data => open,                                                                                    -- (terminated)
			in_empty          => '0',                                                                                     -- (terminated)
			out_empty         => open,                                                                                    -- (terminated)
			in_error          => '0',                                                                                     -- (terminated)
			out_error         => open,                                                                                    -- (terminated)
			in_channel        => '0',                                                                                     -- (terminated)
			out_channel       => open                                                                                     -- (terminated)
		);

	gtp_regif_0_s0_translator_avalon_universal_slave_0_agent : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 58,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 59,
			PKT_TRANS_POSTED          => 60,
			PKT_TRANS_WRITE           => 61,
			PKT_TRANS_READ            => 62,
			PKT_TRANS_LOCK            => 63,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 83,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 68,
			PKT_BYTE_CNT_H            => 67,
			PKT_BYTE_CNT_L            => 65,
			PKT_PROTECTION_H          => 87,
			PKT_PROTECTION_L          => 85,
			PKT_RESPONSE_STATUS_H     => 93,
			PKT_RESPONSE_STATUS_L     => 92,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 94,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                      --       clk_reset.reset
			m0_address              => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_007_src5_ready,                                                       --              cp.ready
			cp_valid                => cmd_xbar_demux_007_src5_valid,                                                       --                .valid
			cp_data                 => cmd_xbar_demux_007_src5_data,                                                        --                .data
			cp_startofpacket        => cmd_xbar_demux_007_src5_startofpacket,                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_007_src5_endofpacket,                                                 --                .endofpacket
			cp_channel              => cmd_xbar_demux_007_src5_channel,                                                     --                .channel
			rf_sink_ready           => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                --     (terminated)
			m0_writeresponserequest => open,                                                                                --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                  --     (terminated)
		);

	gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 95,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_half_clk_clk,                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                      -- clk_reset.reset
			in_data           => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                -- (terminated)
			csr_read          => '0',                                                                                 -- (terminated)
			csr_write         => '0',                                                                                 -- (terminated)
			csr_readdata      => open,                                                                                -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                  -- (terminated)
			almost_full_data  => open,                                                                                -- (terminated)
			almost_empty_data => open,                                                                                -- (terminated)
			in_empty          => '0',                                                                                 -- (terminated)
			out_empty         => open,                                                                                -- (terminated)
			in_error          => '0',                                                                                 -- (terminated)
			out_error         => open,                                                                                -- (terminated)
			in_channel        => '0',                                                                                 -- (terminated)
			out_channel       => open                                                                                 -- (terminated)
		);

	sgdma_tx_csr_translator_avalon_universal_slave_0_agent : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 58,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 59,
			PKT_TRANS_POSTED          => 60,
			PKT_TRANS_WRITE           => 61,
			PKT_TRANS_READ            => 62,
			PKT_TRANS_LOCK            => 63,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 83,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 68,
			PKT_BYTE_CNT_H            => 67,
			PKT_BYTE_CNT_L            => 65,
			PKT_PROTECTION_H          => 87,
			PKT_PROTECTION_L          => 85,
			PKT_RESPONSE_STATUS_H     => 93,
			PKT_RESPONSE_STATUS_L     => 92,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 94,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                          --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                    --       clk_reset.reset
			m0_address              => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_007_src6_ready,                                                     --              cp.ready
			cp_valid                => cmd_xbar_demux_007_src6_valid,                                                     --                .valid
			cp_data                 => cmd_xbar_demux_007_src6_data,                                                      --                .data
			cp_startofpacket        => cmd_xbar_demux_007_src6_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_007_src6_endofpacket,                                               --                .endofpacket
			cp_channel              => cmd_xbar_demux_007_src6_channel,                                                   --                .channel
			rf_sink_ready           => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                --     (terminated)
		);

	sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 95,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_half_clk_clk,                                                          --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			in_data           => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                              -- (terminated)
			csr_read          => '0',                                                                               -- (terminated)
			csr_write         => '0',                                                                               -- (terminated)
			csr_readdata      => open,                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                -- (terminated)
			almost_full_data  => open,                                                                              -- (terminated)
			almost_empty_data => open,                                                                              -- (terminated)
			in_empty          => '0',                                                                               -- (terminated)
			out_empty         => open,                                                                              -- (terminated)
			in_error          => '0',                                                                               -- (terminated)
			out_error         => open,                                                                              -- (terminated)
			in_channel        => '0',                                                                               -- (terminated)
			out_channel       => open                                                                               -- (terminated)
		);

	sgdma_rx_csr_translator_avalon_universal_slave_0_agent : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 76,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 58,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 59,
			PKT_TRANS_POSTED          => 60,
			PKT_TRANS_WRITE           => 61,
			PKT_TRANS_READ            => 62,
			PKT_TRANS_LOCK            => 63,
			PKT_SRC_ID_H              => 80,
			PKT_SRC_ID_L              => 78,
			PKT_DEST_ID_H             => 83,
			PKT_DEST_ID_L             => 81,
			PKT_BURSTWRAP_H           => 68,
			PKT_BURSTWRAP_L           => 68,
			PKT_BYTE_CNT_H            => 67,
			PKT_BYTE_CNT_L            => 65,
			PKT_PROTECTION_H          => 87,
			PKT_PROTECTION_L          => 85,
			PKT_RESPONSE_STATUS_H     => 93,
			PKT_RESPONSE_STATUS_L     => 92,
			PKT_BURST_SIZE_H          => 71,
			PKT_BURST_SIZE_L          => 69,
			ST_CHANNEL_W              => 8,
			ST_DATA_W                 => 94,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                          --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                    --       clk_reset.reset
			m0_address              => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_007_src7_ready,                                                     --              cp.ready
			cp_valid                => cmd_xbar_demux_007_src7_valid,                                                     --                .valid
			cp_data                 => cmd_xbar_demux_007_src7_data,                                                      --                .data
			cp_startofpacket        => cmd_xbar_demux_007_src7_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_007_src7_endofpacket,                                               --                .endofpacket
			cp_channel              => cmd_xbar_demux_007_src7_channel,                                                   --                .channel
			rf_sink_ready           => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                --     (terminated)
		);

	sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 95,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_half_clk_clk,                                                          --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                    -- clk_reset.reset
			in_data           => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                              -- (terminated)
			csr_read          => '0',                                                                               -- (terminated)
			csr_write         => '0',                                                                               -- (terminated)
			csr_readdata      => open,                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                -- (terminated)
			almost_full_data  => open,                                                                              -- (terminated)
			almost_empty_data => open,                                                                              -- (terminated)
			in_empty          => '0',                                                                               -- (terminated)
			out_empty         => open,                                                                              -- (terminated)
			in_error          => '0',                                                                               -- (terminated)
			out_error         => open,                                                                              -- (terminated)
			in_channel        => '0',                                                                               -- (terminated)
			out_channel       => open                                                                               -- (terminated)
		);

	cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent : component sopc_system_cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 88,
			PKT_PROTECTION_L          => 86,
			PKT_BEGIN_BURST           => 81,
			PKT_BURSTWRAP_H           => 73,
			PKT_BURSTWRAP_L           => 73,
			PKT_BURST_SIZE_H          => 76,
			PKT_BURST_SIZE_L          => 74,
			PKT_BURST_TYPE_H          => 78,
			PKT_BURST_TYPE_L          => 77,
			PKT_BYTE_CNT_H            => 72,
			PKT_BYTE_CNT_L            => 70,
			PKT_ADDR_H                => 63,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 64,
			PKT_TRANS_POSTED          => 65,
			PKT_TRANS_WRITE           => 66,
			PKT_TRANS_READ            => 67,
			PKT_TRANS_LOCK            => 68,
			PKT_TRANS_EXCLUSIVE       => 69,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 83,
			PKT_SRC_ID_L              => 83,
			PKT_DEST_ID_H             => 84,
			PKT_DEST_ID_L             => 84,
			PKT_THREAD_ID_H           => 85,
			PKT_THREAD_ID_L           => 85,
			PKT_CACHE_H               => 92,
			PKT_CACHE_L               => 89,
			PKT_DATA_SIDEBAND_H       => 80,
			PKT_DATA_SIDEBAND_L       => 80,
			PKT_QOS_H                 => 82,
			PKT_QOS_L                 => 82,
			PKT_ADDR_SIDEBAND_H       => 79,
			PKT_ADDR_SIDEBAND_L       => 79,
			PKT_RESPONSE_STATUS_H     => 94,
			PKT_RESPONSE_STATUS_L     => 93,
			ST_DATA_W                 => 95,
			ST_CHANNEL_W              => 2,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 1,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                        --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			av_address              => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => limiter_003_rsp_src_valid,                                                       --        rp.valid
			rp_data                 => limiter_003_rsp_src_data,                                                        --          .data
			rp_channel              => limiter_003_rsp_src_channel,                                                     --          .channel
			rp_startofpacket        => limiter_003_rsp_src_startofpacket,                                               --          .startofpacket
			rp_endofpacket          => limiter_003_rsp_src_endofpacket,                                                 --          .endofpacket
			rp_ready                => limiter_003_rsp_src_ready,                                                       --          .ready
			av_response             => open,                                                                            -- (terminated)
			av_writeresponserequest => '0',                                                                             -- (terminated)
			av_writeresponsevalid   => open                                                                             -- (terminated)
		);

	cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent : component sopc_system_cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 63,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 45,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 46,
			PKT_TRANS_POSTED          => 47,
			PKT_TRANS_WRITE           => 48,
			PKT_TRANS_READ            => 49,
			PKT_TRANS_LOCK            => 50,
			PKT_SRC_ID_H              => 65,
			PKT_SRC_ID_L              => 65,
			PKT_DEST_ID_H             => 66,
			PKT_DEST_ID_L             => 66,
			PKT_BURSTWRAP_H           => 55,
			PKT_BURSTWRAP_L           => 55,
			PKT_BYTE_CNT_H            => 54,
			PKT_BYTE_CNT_L            => 52,
			PKT_PROTECTION_H          => 70,
			PKT_PROTECTION_L          => 68,
			PKT_RESPONSE_STATUS_H     => 76,
			PKT_RESPONSE_STATUS_L     => 75,
			PKT_BURST_SIZE_H          => 58,
			PKT_BURST_SIZE_L          => 56,
			ST_CHANNEL_W              => 2,
			ST_DATA_W                 => 77,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                                              --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                        --       clk_reset.reset
			m0_address              => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_source0_ready,                                                                           --              cp.ready
			cp_valid                => burst_adapter_source0_valid,                                                                           --                .valid
			cp_data                 => burst_adapter_source0_data,                                                                            --                .data
			cp_startofpacket        => burst_adapter_source0_startofpacket,                                                                   --                .startofpacket
			cp_endofpacket          => burst_adapter_source0_endofpacket,                                                                     --                .endofpacket
			cp_channel              => burst_adapter_source0_channel,                                                                         --                .channel
			rf_sink_ready           => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                  --     (terminated)
			m0_writeresponserequest => open,                                                                                                  --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                    --     (terminated)
		);

	cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 78,
			FIFO_DEPTH          => 4,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_half_clk_clk,                                                                              --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                        -- clk_reset.reset
			in_data           => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                  -- (terminated)
			csr_read          => '0',                                                                                                   -- (terminated)
			csr_write         => '0',                                                                                                   -- (terminated)
			csr_readdata      => open,                                                                                                  -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                    -- (terminated)
			almost_full_data  => open,                                                                                                  -- (terminated)
			almost_empty_data => open,                                                                                                  -- (terminated)
			in_empty          => '0',                                                                                                   -- (terminated)
			out_empty         => open,                                                                                                  -- (terminated)
			in_error          => '0',                                                                                                   -- (terminated)
			out_error         => open,                                                                                                  -- (terminated)
			in_channel        => '0',                                                                                                   -- (terminated)
			out_channel       => open                                                                                                   -- (terminated)
		);

	cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo : component sopc_system_cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 18,
			FIFO_DEPTH          => 4,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_half_clk_clk,                                                                        --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                  -- clk_reset.reset
			in_data           => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                                            -- (terminated)
			csr_read          => '0',                                                                                             -- (terminated)
			csr_write         => '0',                                                                                             -- (terminated)
			csr_readdata      => open,                                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                              -- (terminated)
			almost_full_data  => open,                                                                                            -- (terminated)
			almost_empty_data => open,                                                                                            -- (terminated)
			in_startofpacket  => '0',                                                                                             -- (terminated)
			in_endofpacket    => '0',                                                                                             -- (terminated)
			out_startofpacket => open,                                                                                            -- (terminated)
			out_endofpacket   => open,                                                                                            -- (terminated)
			in_empty          => '0',                                                                                             -- (terminated)
			out_empty         => open,                                                                                            -- (terminated)
			in_error          => '0',                                                                                             -- (terminated)
			out_error         => open,                                                                                            -- (terminated)
			in_channel        => '0',                                                                                             -- (terminated)
			out_channel       => open                                                                                             -- (terminated)
		);

	cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent : component sopc_system_cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 63,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 45,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 46,
			PKT_TRANS_POSTED          => 47,
			PKT_TRANS_WRITE           => 48,
			PKT_TRANS_READ            => 49,
			PKT_TRANS_LOCK            => 50,
			PKT_SRC_ID_H              => 65,
			PKT_SRC_ID_L              => 65,
			PKT_DEST_ID_H             => 66,
			PKT_DEST_ID_L             => 66,
			PKT_BURSTWRAP_H           => 55,
			PKT_BURSTWRAP_L           => 55,
			PKT_BYTE_CNT_H            => 54,
			PKT_BYTE_CNT_L            => 52,
			PKT_PROTECTION_H          => 70,
			PKT_PROTECTION_L          => 68,
			PKT_RESPONSE_STATUS_H     => 76,
			PKT_RESPONSE_STATUS_L     => 75,
			PKT_BURST_SIZE_H          => 58,
			PKT_BURST_SIZE_L          => 56,
			ST_CHANNEL_W              => 2,
			ST_DATA_W                 => 77,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                   --       clk_reset.reset
			m0_address              => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_001_source0_ready,                                                                  --              cp.ready
			cp_valid                => burst_adapter_001_source0_valid,                                                                  --                .valid
			cp_data                 => burst_adapter_001_source0_data,                                                                   --                .data
			cp_startofpacket        => burst_adapter_001_source0_startofpacket,                                                          --                .startofpacket
			cp_endofpacket          => burst_adapter_001_source0_endofpacket,                                                            --                .endofpacket
			cp_channel              => burst_adapter_001_source0_channel,                                                                --                .channel
			rf_sink_ready           => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                               --     (terminated)
		);

	cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 78,
			FIFO_DEPTH          => 4,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_half_clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                   -- clk_reset.reset
			in_data           => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                             -- (terminated)
			csr_read          => '0',                                                                                              -- (terminated)
			csr_write         => '0',                                                                                              -- (terminated)
			csr_readdata      => open,                                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                               -- (terminated)
			almost_full_data  => open,                                                                                             -- (terminated)
			almost_empty_data => open,                                                                                             -- (terminated)
			in_empty          => '0',                                                                                              -- (terminated)
			out_empty         => open,                                                                                             -- (terminated)
			in_error          => '0',                                                                                              -- (terminated)
			out_error         => open,                                                                                             -- (terminated)
			in_channel        => '0',                                                                                              -- (terminated)
			out_channel       => open                                                                                              -- (terminated)
		);

	cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo : component sopc_system_cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 18,
			FIFO_DEPTH          => 4,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_half_clk_clk,                                                                   --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                             -- clk_reset.reset
			in_data           => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                                       -- (terminated)
			csr_read          => '0',                                                                                        -- (terminated)
			csr_write         => '0',                                                                                        -- (terminated)
			csr_readdata      => open,                                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                         -- (terminated)
			almost_full_data  => open,                                                                                       -- (terminated)
			almost_empty_data => open,                                                                                       -- (terminated)
			in_startofpacket  => '0',                                                                                        -- (terminated)
			in_endofpacket    => '0',                                                                                        -- (terminated)
			out_startofpacket => open,                                                                                       -- (terminated)
			out_endofpacket   => open,                                                                                       -- (terminated)
			in_empty          => '0',                                                                                        -- (terminated)
			out_empty         => open,                                                                                       -- (terminated)
			in_error          => '0',                                                                                        -- (terminated)
			out_error         => open,                                                                                       -- (terminated)
			in_channel        => '0',                                                                                        -- (terminated)
			out_channel       => open                                                                                        -- (terminated)
		);

	sgdma_tx_m_read_translator_avalon_universal_master_0_agent : component sopc_system_sgdma_tx_m_read_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 92,
			PKT_PROTECTION_L          => 90,
			PKT_BEGIN_BURST           => 85,
			PKT_BURSTWRAP_H           => 77,
			PKT_BURSTWRAP_L           => 77,
			PKT_BURST_SIZE_H          => 80,
			PKT_BURST_SIZE_L          => 78,
			PKT_BURST_TYPE_H          => 82,
			PKT_BURST_TYPE_L          => 81,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 87,
			PKT_DEST_ID_H             => 88,
			PKT_DEST_ID_L             => 88,
			PKT_THREAD_ID_H           => 89,
			PKT_THREAD_ID_L           => 89,
			PKT_CACHE_H               => 96,
			PKT_CACHE_L               => 93,
			PKT_DATA_SIDEBAND_H       => 84,
			PKT_DATA_SIDEBAND_L       => 84,
			PKT_QOS_H                 => 86,
			PKT_QOS_L                 => 86,
			PKT_ADDR_SIDEBAND_H       => 83,
			PKT_ADDR_SIDEBAND_L       => 83,
			PKT_RESPONSE_STATUS_H     => 98,
			PKT_RESPONSE_STATUS_L     => 97,
			ST_DATA_W                 => 99,
			ST_CHANNEL_W              => 2,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 1,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                    --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			av_address              => sgdma_tx_m_read_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => sgdma_tx_m_read_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => sgdma_tx_m_read_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => sgdma_tx_m_read_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => sgdma_tx_m_read_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => sgdma_tx_m_read_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => sgdma_tx_m_read_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => sgdma_tx_m_read_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => sgdma_tx_m_read_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => sgdma_tx_m_read_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => sgdma_tx_m_read_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_demux_015_src0_valid,                                               --        rp.valid
			rp_data                 => rsp_xbar_demux_015_src0_data,                                                --          .data
			rp_channel              => rsp_xbar_demux_015_src0_channel,                                             --          .channel
			rp_startofpacket        => rsp_xbar_demux_015_src0_startofpacket,                                       --          .startofpacket
			rp_endofpacket          => rsp_xbar_demux_015_src0_endofpacket,                                         --          .endofpacket
			rp_ready                => rsp_xbar_demux_015_src0_ready,                                               --          .ready
			av_response             => open,                                                                        -- (terminated)
			av_writeresponserequest => '0',                                                                         -- (terminated)
			av_writeresponsevalid   => open                                                                         -- (terminated)
		);

	sgdma_rx_m_write_translator_avalon_universal_master_0_agent : component sopc_system_sgdma_tx_m_read_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 92,
			PKT_PROTECTION_L          => 90,
			PKT_BEGIN_BURST           => 85,
			PKT_BURSTWRAP_H           => 77,
			PKT_BURSTWRAP_L           => 77,
			PKT_BURST_SIZE_H          => 80,
			PKT_BURST_SIZE_L          => 78,
			PKT_BURST_TYPE_H          => 82,
			PKT_BURST_TYPE_L          => 81,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_TRANS_EXCLUSIVE       => 73,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 87,
			PKT_DEST_ID_H             => 88,
			PKT_DEST_ID_L             => 88,
			PKT_THREAD_ID_H           => 89,
			PKT_THREAD_ID_L           => 89,
			PKT_CACHE_H               => 96,
			PKT_CACHE_L               => 93,
			PKT_DATA_SIDEBAND_H       => 84,
			PKT_DATA_SIDEBAND_L       => 84,
			PKT_QOS_H                 => 86,
			PKT_QOS_L                 => 86,
			PKT_ADDR_SIDEBAND_H       => 83,
			PKT_ADDR_SIDEBAND_L       => 83,
			PKT_RESPONSE_STATUS_H     => 98,
			PKT_RESPONSE_STATUS_L     => 97,
			ST_DATA_W                 => 99,
			ST_CHANNEL_W              => 2,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 1,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                     --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                               -- clk_reset.reset
			av_address              => sgdma_rx_m_write_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => sgdma_rx_m_write_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => sgdma_rx_m_write_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => sgdma_rx_m_write_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => sgdma_rx_m_write_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => sgdma_rx_m_write_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => sgdma_rx_m_write_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => sgdma_rx_m_write_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => sgdma_rx_m_write_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => sgdma_rx_m_write_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => sgdma_rx_m_write_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_demux_015_src1_valid,                                                --        rp.valid
			rp_data                 => rsp_xbar_demux_015_src1_data,                                                 --          .data
			rp_channel              => rsp_xbar_demux_015_src1_channel,                                              --          .channel
			rp_startofpacket        => rsp_xbar_demux_015_src1_startofpacket,                                        --          .startofpacket
			rp_endofpacket          => rsp_xbar_demux_015_src1_endofpacket,                                          --          .endofpacket
			rp_ready                => rsp_xbar_demux_015_src1_ready,                                                --          .ready
			av_response             => open,                                                                         -- (terminated)
			av_writeresponserequest => '0',                                                                          -- (terminated)
			av_writeresponsevalid   => open                                                                          -- (terminated)
		);

	tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent : component sopc_system_tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 85,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 67,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 68,
			PKT_TRANS_POSTED          => 69,
			PKT_TRANS_WRITE           => 70,
			PKT_TRANS_READ            => 71,
			PKT_TRANS_LOCK            => 72,
			PKT_SRC_ID_H              => 87,
			PKT_SRC_ID_L              => 87,
			PKT_DEST_ID_H             => 88,
			PKT_DEST_ID_L             => 88,
			PKT_BURSTWRAP_H           => 77,
			PKT_BURSTWRAP_L           => 77,
			PKT_BYTE_CNT_H            => 76,
			PKT_BYTE_CNT_L            => 74,
			PKT_PROTECTION_H          => 92,
			PKT_PROTECTION_L          => 90,
			PKT_RESPONSE_STATUS_H     => 98,
			PKT_RESPONSE_STATUS_L     => 97,
			PKT_BURST_SIZE_H          => 80,
			PKT_BURST_SIZE_L          => 78,
			ST_CHANNEL_W              => 2,
			ST_DATA_W                 => 99,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_half_clk_clk,                                                                     --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                               --       clk_reset.reset
			m0_address              => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_015_src_ready,                                                                   --              cp.ready
			cp_valid                => cmd_xbar_mux_015_src_valid,                                                                   --                .valid
			cp_data                 => cmd_xbar_mux_015_src_data,                                                                    --                .data
			cp_startofpacket        => cmd_xbar_mux_015_src_startofpacket,                                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_015_src_endofpacket,                                                             --                .endofpacket
			cp_channel              => cmd_xbar_mux_015_src_channel,                                                                 --                .channel
			rf_sink_ready           => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                         --     (terminated)
			m0_writeresponserequest => open,                                                                                         --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                           --     (terminated)
		);

	tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 100,
			FIFO_DEPTH          => 9,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_half_clk_clk,                                                                     --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                               -- clk_reset.reset
			in_data           => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                         -- (terminated)
			csr_read          => '0',                                                                                          -- (terminated)
			csr_write         => '0',                                                                                          -- (terminated)
			csr_readdata      => open,                                                                                         -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                           -- (terminated)
			almost_full_data  => open,                                                                                         -- (terminated)
			almost_empty_data => open,                                                                                         -- (terminated)
			in_empty          => '0',                                                                                          -- (terminated)
			out_empty         => open,                                                                                         -- (terminated)
			in_error          => '0',                                                                                          -- (terminated)
			out_error         => open,                                                                                         -- (terminated)
			in_channel        => '0',                                                                                          -- (terminated)
			out_channel       => open                                                                                          -- (terminated)
		);

	tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent : component sopc_system_tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 90,
			PKT_PROTECTION_L          => 88,
			PKT_BEGIN_BURST           => 83,
			PKT_BURSTWRAP_H           => 75,
			PKT_BURSTWRAP_L           => 75,
			PKT_BURST_SIZE_H          => 78,
			PKT_BURST_SIZE_L          => 76,
			PKT_BURST_TYPE_H          => 80,
			PKT_BURST_TYPE_L          => 79,
			PKT_BYTE_CNT_H            => 74,
			PKT_BYTE_CNT_L            => 69,
			PKT_ADDR_H                => 62,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 63,
			PKT_TRANS_POSTED          => 64,
			PKT_TRANS_WRITE           => 65,
			PKT_TRANS_READ            => 66,
			PKT_TRANS_LOCK            => 67,
			PKT_TRANS_EXCLUSIVE       => 68,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 85,
			PKT_DEST_ID_H             => 86,
			PKT_DEST_ID_L             => 86,
			PKT_THREAD_ID_H           => 87,
			PKT_THREAD_ID_L           => 87,
			PKT_CACHE_H               => 94,
			PKT_CACHE_L               => 91,
			PKT_DATA_SIDEBAND_H       => 82,
			PKT_DATA_SIDEBAND_L       => 82,
			PKT_QOS_H                 => 84,
			PKT_QOS_L                 => 84,
			PKT_ADDR_SIDEBAND_H       => 81,
			PKT_ADDR_SIDEBAND_L       => 81,
			PKT_RESPONSE_STATUS_H     => 96,
			PKT_RESPONSE_STATUS_L     => 95,
			ST_DATA_W                 => 97,
			ST_CHANNEL_W              => 2,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 1,
			ID                        => 1,
			BURSTWRAP_VALUE           => 1,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_clk_clk,                                                                 --       clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                  -- clk_reset.reset
			av_address              => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_demux_016_src0_valid,                                                       --        rp.valid
			rp_data                 => rsp_xbar_demux_016_src0_data,                                                        --          .data
			rp_channel              => rsp_xbar_demux_016_src0_channel,                                                     --          .channel
			rp_startofpacket        => rsp_xbar_demux_016_src0_startofpacket,                                               --          .startofpacket
			rp_endofpacket          => rsp_xbar_demux_016_src0_endofpacket,                                                 --          .endofpacket
			rp_ready                => rsp_xbar_demux_016_src0_ready,                                                       --          .ready
			av_response             => open,                                                                                -- (terminated)
			av_writeresponserequest => '0',                                                                                 -- (terminated)
			av_writeresponsevalid   => open                                                                                 -- (terminated)
		);

	cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent : component sopc_system_tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent
		generic map (
			PKT_PROTECTION_H          => 90,
			PKT_PROTECTION_L          => 88,
			PKT_BEGIN_BURST           => 83,
			PKT_BURSTWRAP_H           => 75,
			PKT_BURSTWRAP_L           => 75,
			PKT_BURST_SIZE_H          => 78,
			PKT_BURST_SIZE_L          => 76,
			PKT_BURST_TYPE_H          => 80,
			PKT_BURST_TYPE_L          => 79,
			PKT_BYTE_CNT_H            => 74,
			PKT_BYTE_CNT_L            => 69,
			PKT_ADDR_H                => 62,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 63,
			PKT_TRANS_POSTED          => 64,
			PKT_TRANS_WRITE           => 65,
			PKT_TRANS_READ            => 66,
			PKT_TRANS_LOCK            => 67,
			PKT_TRANS_EXCLUSIVE       => 68,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 85,
			PKT_SRC_ID_L              => 85,
			PKT_DEST_ID_H             => 86,
			PKT_DEST_ID_L             => 86,
			PKT_THREAD_ID_H           => 87,
			PKT_THREAD_ID_L           => 87,
			PKT_CACHE_H               => 94,
			PKT_CACHE_L               => 91,
			PKT_DATA_SIDEBAND_H       => 82,
			PKT_DATA_SIDEBAND_L       => 82,
			PKT_QOS_H                 => 84,
			PKT_QOS_L                 => 84,
			PKT_ADDR_SIDEBAND_H       => 81,
			PKT_ADDR_SIDEBAND_L       => 81,
			PKT_RESPONSE_STATUS_H     => 96,
			PKT_RESPONSE_STATUS_L     => 95,
			ST_DATA_W                 => 97,
			ST_CHANNEL_W              => 2,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 1,
			ID                        => 0,
			BURSTWRAP_VALUE           => 1,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_clk_clk,                                                            --       clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                             -- clk_reset.reset
			av_address              => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_demux_016_src1_valid,                                                  --        rp.valid
			rp_data                 => rsp_xbar_demux_016_src1_data,                                                   --          .data
			rp_channel              => rsp_xbar_demux_016_src1_channel,                                                --          .channel
			rp_startofpacket        => rsp_xbar_demux_016_src1_startofpacket,                                          --          .startofpacket
			rp_endofpacket          => rsp_xbar_demux_016_src1_endofpacket,                                            --          .endofpacket
			rp_ready                => rsp_xbar_demux_016_src1_ready,                                                  --          .ready
			av_response             => open,                                                                           -- (terminated)
			av_writeresponserequest => '0',                                                                            -- (terminated)
			av_writeresponsevalid   => open                                                                            -- (terminated)
		);

	sdram_0_avl_translator_avalon_universal_slave_0_agent : component sopc_system_sdram_0_avl_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 63,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 119,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 71,
			PKT_BYTEEN_L              => 64,
			PKT_ADDR_H                => 98,
			PKT_ADDR_L                => 72,
			PKT_TRANS_COMPRESSED_READ => 99,
			PKT_TRANS_POSTED          => 100,
			PKT_TRANS_WRITE           => 101,
			PKT_TRANS_READ            => 102,
			PKT_TRANS_LOCK            => 103,
			PKT_SRC_ID_H              => 121,
			PKT_SRC_ID_L              => 121,
			PKT_DEST_ID_H             => 122,
			PKT_DEST_ID_L             => 122,
			PKT_BURSTWRAP_H           => 111,
			PKT_BURSTWRAP_L           => 111,
			PKT_BYTE_CNT_H            => 110,
			PKT_BYTE_CNT_L            => 105,
			PKT_PROTECTION_H          => 126,
			PKT_PROTECTION_L          => 124,
			PKT_RESPONSE_STATUS_H     => 132,
			PKT_RESPONSE_STATUS_L     => 131,
			PKT_BURST_SIZE_H          => 114,
			PKT_BURST_SIZE_L          => 112,
			ST_CHANNEL_W              => 2,
			ST_DATA_W                 => 133,
			AVS_BURSTCOUNT_W          => 6,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => sdram_0_afi_clk_clk,                                                              --             clk.clk
			reset                   => rst_controller_004_reset_out_reset,                                               --       clk_reset.reset
			m0_address              => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sdram_0_avl_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sdram_0_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sdram_0_avl_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sdram_0_avl_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sdram_0_avl_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sdram_0_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => width_adapter_004_src_ready,                                                      --              cp.ready
			cp_valid                => width_adapter_004_src_valid,                                                      --                .valid
			cp_data                 => width_adapter_004_src_data,                                                       --                .data
			cp_startofpacket        => width_adapter_004_src_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => width_adapter_004_src_endofpacket,                                                --                .endofpacket
			cp_channel              => width_adapter_004_src_channel,                                                    --                .channel
			rf_sink_ready           => sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sdram_0_avl_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sdram_0_avl_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sdram_0_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sdram_0_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sdram_0_avl_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sdram_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sdram_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sdram_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sdram_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sdram_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sdram_0_avl_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                               --     (terminated)
		);

	sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo : component sopc_system_sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 134,
			FIFO_DEPTH          => 33,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => sdram_0_afi_clk_clk,                                                              --       clk.clk
			reset             => rst_controller_004_reset_out_reset,                                               -- clk_reset.reset
			in_data           => sdram_0_avl_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sdram_0_avl_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sdram_0_avl_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sdram_0_avl_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sdram_0_avl_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sdram_0_avl_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                             -- (terminated)
			csr_read          => '0',                                                                              -- (terminated)
			csr_write         => '0',                                                                              -- (terminated)
			csr_readdata      => open,                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                               -- (terminated)
			almost_full_data  => open,                                                                             -- (terminated)
			almost_empty_data => open,                                                                             -- (terminated)
			in_empty          => '0',                                                                              -- (terminated)
			out_empty         => open,                                                                             -- (terminated)
			in_error          => '0',                                                                              -- (terminated)
			out_error         => open,                                                                             -- (terminated)
			in_channel        => '0',                                                                              -- (terminated)
			out_channel       => open                                                                              -- (terminated)
		);

	addr_router : component sopc_system_addr_router
		port map (
			sink_ready         => linux_cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => linux_cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => linux_cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => linux_cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => linux_cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_clk_clk,                                                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                             --       src.ready
			src_valid          => addr_router_src_valid,                                                             --          .valid
			src_data           => addr_router_src_data,                                                              --          .data
			src_channel        => addr_router_src_channel,                                                           --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                     --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                        --          .endofpacket
		);

	addr_router_001 : component sopc_system_addr_router_001
		port map (
			sink_ready         => linux_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => linux_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => linux_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => linux_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => linux_cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_clk_clk,                                                                      --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                       -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                                --       src.ready
			src_valid          => addr_router_001_src_valid,                                                                --          .valid
			src_data           => addr_router_001_src_data,                                                                 --          .data
			src_channel        => addr_router_001_src_channel,                                                              --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                                           --          .endofpacket
		);

	id_router : component sopc_system_id_router
		port map (
			sink_ready         => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => linux_cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_clk_clk,                                                                    --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                                    --       src.ready
			src_valid          => id_router_src_valid,                                                                    --          .valid
			src_data           => id_router_src_data,                                                                     --          .data
			src_channel        => id_router_src_channel,                                                                  --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                            --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                               --          .endofpacket
		);

	id_router_001 : component sopc_system_id_router
		port map (
			sink_ready         => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_to_flash_ccb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_clk_clk,                                                            --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                             -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                                        --       src.ready
			src_valid          => id_router_001_src_valid,                                                        --          .valid
			src_data           => id_router_001_src_data,                                                         --          .data
			src_channel        => id_router_001_src_channel,                                                      --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                                --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                                   --          .endofpacket
		);

	id_router_002 : component sopc_system_id_router_002
		port map (
			sink_ready         => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_to_peripherals_ccb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_clk_clk,                                                                  --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                   -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                              --       src.ready
			src_valid          => id_router_002_src_valid,                                                              --          .valid
			src_data           => id_router_002_src_data,                                                               --          .data
			src_channel        => id_router_002_src_channel,                                                            --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                         --          .endofpacket
		);

	id_router_003 : component sopc_system_id_router
		port map (
			sink_ready         => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_to_sdram_pb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_clk_clk,                                                           --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                            -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                       --       src.ready
			src_valid          => id_router_003_src_valid,                                                       --          .valid
			src_data           => id_router_003_src_data,                                                        --          .data
			src_channel        => id_router_003_src_channel,                                                     --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                               --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                                  --          .endofpacket
		);

	addr_router_002 : component sopc_system_addr_router_002
		port map (
			sink_ready         => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => sgdma_tx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			src_ready          => addr_router_002_src_ready,                                                             --       src.ready
			src_valid          => addr_router_002_src_valid,                                                             --          .valid
			src_data           => addr_router_002_src_data,                                                              --          .data
			src_channel        => addr_router_002_src_channel,                                                           --          .channel
			src_startofpacket  => addr_router_002_src_startofpacket,                                                     --          .startofpacket
			src_endofpacket    => addr_router_002_src_endofpacket                                                        --          .endofpacket
		);

	addr_router_003 : component sopc_system_addr_router_002
		port map (
			sink_ready         => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => sgdma_rx_descriptor_write_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			src_ready          => addr_router_003_src_ready,                                                             --       src.ready
			src_valid          => addr_router_003_src_valid,                                                             --          .valid
			src_data           => addr_router_003_src_data,                                                              --          .data
			src_channel        => addr_router_003_src_channel,                                                           --          .channel
			src_startofpacket  => addr_router_003_src_startofpacket,                                                     --          .startofpacket
			src_endofpacket    => addr_router_003_src_endofpacket                                                        --          .endofpacket
		);

	addr_router_004 : component sopc_system_addr_router_002
		port map (
			sink_ready         => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => sgdma_rx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                             --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			src_ready          => addr_router_004_src_ready,                                                            --       src.ready
			src_valid          => addr_router_004_src_valid,                                                            --          .valid
			src_data           => addr_router_004_src_data,                                                             --          .data
			src_channel        => addr_router_004_src_channel,                                                          --          .channel
			src_startofpacket  => addr_router_004_src_startofpacket,                                                    --          .startofpacket
			src_endofpacket    => addr_router_004_src_endofpacket                                                       --          .endofpacket
		);

	addr_router_005 : component sopc_system_addr_router_002
		port map (
			sink_ready         => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => sgdma_tx_descriptor_read_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                             --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			src_ready          => addr_router_005_src_ready,                                                            --       src.ready
			src_valid          => addr_router_005_src_valid,                                                            --          .valid
			src_data           => addr_router_005_src_data,                                                             --          .data
			src_channel        => addr_router_005_src_channel,                                                          --          .channel
			src_startofpacket  => addr_router_005_src_startofpacket,                                                    --          .startofpacket
			src_endofpacket    => addr_router_005_src_endofpacket                                                       --          .endofpacket
		);

	id_router_004 : component sopc_system_id_router_004
		port map (
			sink_ready         => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => dma_to_descriptor_mem_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                      -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                                             --       src.ready
			src_valid          => id_router_004_src_valid,                                                             --          .valid
			src_data           => id_router_004_src_data,                                                              --          .data
			src_channel        => id_router_004_src_channel,                                                           --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                                     --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                                        --          .endofpacket
		);

	addr_router_006 : component sopc_system_addr_router_006
		port map (
			sink_ready         => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => dma_to_descriptor_mem_m0_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                             --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			src_ready          => addr_router_006_src_ready,                                                            --       src.ready
			src_valid          => addr_router_006_src_valid,                                                            --          .valid
			src_data           => addr_router_006_src_data,                                                             --          .data
			src_channel        => addr_router_006_src_channel,                                                          --          .channel
			src_startofpacket  => addr_router_006_src_startofpacket,                                                    --          .startofpacket
			src_endofpacket    => addr_router_006_src_endofpacket                                                       --          .endofpacket
		);

	addr_router_007 : component sopc_system_addr_router_007
		port map (
			sink_ready         => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_to_peripherals_ccb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			src_ready          => addr_router_007_src_ready,                                                             --       src.ready
			src_valid          => addr_router_007_src_valid,                                                             --          .valid
			src_data           => addr_router_007_src_data,                                                              --          .data
			src_channel        => addr_router_007_src_channel,                                                           --          .channel
			src_startofpacket  => addr_router_007_src_startofpacket,                                                     --          .startofpacket
			src_endofpacket    => addr_router_007_src_endofpacket                                                        --          .endofpacket
		);

	id_router_005 : component sopc_system_id_router_005
		port map (
			sink_ready         => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => descriptor_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                        --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                                         --       src.ready
			src_valid          => id_router_005_src_valid,                                                         --          .valid
			src_data           => id_router_005_src_data,                                                          --          .data
			src_channel        => id_router_005_src_channel,                                                       --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                                 --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                                    --          .endofpacket
		);

	id_router_006 : component sopc_system_id_router_006
		port map (
			sink_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                                                --       src.ready
			src_valid          => id_router_006_src_valid,                                                                --          .valid
			src_data           => id_router_006_src_data,                                                                 --          .data
			src_channel        => id_router_006_src_channel,                                                              --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                                           --          .endofpacket
		);

	id_router_007 : component sopc_system_id_router_006
		port map (
			sink_ready         => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => tse_mac_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                        --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                                         --       src.ready
			src_valid          => id_router_007_src_valid,                                                         --          .valid
			src_data           => id_router_007_src_data,                                                          --          .data
			src_channel        => id_router_007_src_channel,                                                       --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                                 --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                                    --          .endofpacket
		);

	id_router_008 : component sopc_system_id_router_006
		port map (
			sink_ready         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                       --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			src_ready          => id_router_008_src_ready,                                                        --       src.ready
			src_valid          => id_router_008_src_valid,                                                        --          .valid
			src_data           => id_router_008_src_data,                                                         --          .data
			src_channel        => id_router_008_src_channel,                                                      --          .channel
			src_startofpacket  => id_router_008_src_startofpacket,                                                --          .startofpacket
			src_endofpacket    => id_router_008_src_endofpacket                                                   --          .endofpacket
		);

	id_router_009 : component sopc_system_id_router_006
		port map (
			sink_ready         => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => linux_timer_1ms_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                      --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                -- clk_reset.reset
			src_ready          => id_router_009_src_ready,                                                       --       src.ready
			src_valid          => id_router_009_src_valid,                                                       --          .valid
			src_data           => id_router_009_src_data,                                                        --          .data
			src_channel        => id_router_009_src_channel,                                                     --          .channel
			src_startofpacket  => id_router_009_src_startofpacket,                                               --          .startofpacket
			src_endofpacket    => id_router_009_src_endofpacket                                                  --          .endofpacket
		);

	id_router_010 : component sopc_system_id_router_006
		port map (
			sink_ready         => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => gtp_regif_0_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                            -- clk_reset.reset
			src_ready          => id_router_010_src_ready,                                                   --       src.ready
			src_valid          => id_router_010_src_valid,                                                   --          .valid
			src_data           => id_router_010_src_data,                                                    --          .data
			src_channel        => id_router_010_src_channel,                                                 --          .channel
			src_startofpacket  => id_router_010_src_startofpacket,                                           --          .startofpacket
			src_endofpacket    => id_router_010_src_endofpacket                                              --          .endofpacket
		);

	id_router_011 : component sopc_system_id_router_006
		port map (
			sink_ready         => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sgdma_tx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                --       clk.clk
			reset              => rst_controller_reset_out_reset,                                          -- clk_reset.reset
			src_ready          => id_router_011_src_ready,                                                 --       src.ready
			src_valid          => id_router_011_src_valid,                                                 --          .valid
			src_data           => id_router_011_src_data,                                                  --          .data
			src_channel        => id_router_011_src_channel,                                               --          .channel
			src_startofpacket  => id_router_011_src_startofpacket,                                         --          .startofpacket
			src_endofpacket    => id_router_011_src_endofpacket                                            --          .endofpacket
		);

	id_router_012 : component sopc_system_id_router_006
		port map (
			sink_ready         => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sgdma_rx_csr_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                --       clk.clk
			reset              => rst_controller_reset_out_reset,                                          -- clk_reset.reset
			src_ready          => id_router_012_src_ready,                                                 --       src.ready
			src_valid          => id_router_012_src_valid,                                                 --          .valid
			src_data           => id_router_012_src_data,                                                  --          .data
			src_channel        => id_router_012_src_channel,                                               --          .channel
			src_startofpacket  => id_router_012_src_startofpacket,                                         --          .startofpacket
			src_endofpacket    => id_router_012_src_endofpacket                                            --          .endofpacket
		);

	addr_router_008 : component sopc_system_addr_router_008
		port map (
			sink_ready         => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_to_flash_ccb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                        --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			src_ready          => addr_router_008_src_ready,                                                       --       src.ready
			src_valid          => addr_router_008_src_valid,                                                       --          .valid
			src_data           => addr_router_008_src_data,                                                        --          .data
			src_channel        => addr_router_008_src_channel,                                                     --          .channel
			src_startofpacket  => addr_router_008_src_startofpacket,                                               --          .startofpacket
			src_endofpacket    => addr_router_008_src_endofpacket                                                  --          .endofpacket
		);

	id_router_013 : component sopc_system_id_router_013
		port map (
			sink_ready         => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => cfi_flash_ts_controller_fpga_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                                    --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                              -- clk_reset.reset
			src_ready          => id_router_013_src_ready,                                                                     --       src.ready
			src_valid          => id_router_013_src_valid,                                                                     --          .valid
			src_data           => id_router_013_src_data,                                                                      --          .data
			src_channel        => id_router_013_src_channel,                                                                   --          .channel
			src_startofpacket  => id_router_013_src_startofpacket,                                                             --          .startofpacket
			src_endofpacket    => id_router_013_src_endofpacket                                                                --          .endofpacket
		);

	id_router_014 : component sopc_system_id_router_013
		port map (
			sink_ready         => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => cfi_flash_ts_controller_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			src_ready          => id_router_014_src_ready,                                                                --       src.ready
			src_valid          => id_router_014_src_valid,                                                                --          .valid
			src_data           => id_router_014_src_data,                                                                 --          .data
			src_channel        => id_router_014_src_channel,                                                              --          .channel
			src_startofpacket  => id_router_014_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => id_router_014_src_endofpacket                                                           --          .endofpacket
		);

	addr_router_009 : component sopc_system_addr_router_009
		port map (
			sink_ready         => sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => sgdma_tx_m_read_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                    --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => addr_router_009_src_ready,                                                   --       src.ready
			src_valid          => addr_router_009_src_valid,                                                   --          .valid
			src_data           => addr_router_009_src_data,                                                    --          .data
			src_channel        => addr_router_009_src_channel,                                                 --          .channel
			src_startofpacket  => addr_router_009_src_startofpacket,                                           --          .startofpacket
			src_endofpacket    => addr_router_009_src_endofpacket                                              --          .endofpacket
		);

	addr_router_010 : component sopc_system_addr_router_009
		port map (
			sink_ready         => sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => sgdma_rx_m_write_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                               -- clk_reset.reset
			src_ready          => addr_router_010_src_ready,                                                    --       src.ready
			src_valid          => addr_router_010_src_valid,                                                    --          .valid
			src_data           => addr_router_010_src_data,                                                     --          .data
			src_channel        => addr_router_010_src_channel,                                                  --          .channel
			src_startofpacket  => addr_router_010_src_startofpacket,                                            --          .startofpacket
			src_endofpacket    => addr_router_010_src_endofpacket                                               --          .endofpacket
		);

	id_router_015 : component sopc_system_id_router_015
		port map (
			sink_ready         => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => tse_dma_to_sdram_ccb_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_half_clk_clk,                                                           --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => id_router_015_src_ready,                                                            --       src.ready
			src_valid          => id_router_015_src_valid,                                                            --          .valid
			src_data           => id_router_015_src_data,                                                             --          .data
			src_channel        => id_router_015_src_channel,                                                          --          .channel
			src_startofpacket  => id_router_015_src_startofpacket,                                                    --          .startofpacket
			src_endofpacket    => id_router_015_src_endofpacket                                                       --          .endofpacket
		);

	addr_router_011 : component sopc_system_addr_router_011
		port map (
			sink_ready         => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => tse_dma_to_sdram_ccb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_clk_clk,                                                                 --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                  -- clk_reset.reset
			src_ready          => addr_router_011_src_ready,                                                           --       src.ready
			src_valid          => addr_router_011_src_valid,                                                           --          .valid
			src_data           => addr_router_011_src_data,                                                            --          .data
			src_channel        => addr_router_011_src_channel,                                                         --          .channel
			src_startofpacket  => addr_router_011_src_startofpacket,                                                   --          .startofpacket
			src_endofpacket    => addr_router_011_src_endofpacket                                                      --          .endofpacket
		);

	addr_router_012 : component sopc_system_addr_router_011
		port map (
			sink_ready         => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_to_sdram_pb_m0_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_clk_clk,                                                            --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                             -- clk_reset.reset
			src_ready          => addr_router_012_src_ready,                                                      --       src.ready
			src_valid          => addr_router_012_src_valid,                                                      --          .valid
			src_data           => addr_router_012_src_data,                                                       --          .data
			src_channel        => addr_router_012_src_channel,                                                    --          .channel
			src_startofpacket  => addr_router_012_src_startofpacket,                                              --          .startofpacket
			src_endofpacket    => addr_router_012_src_endofpacket                                                 --          .endofpacket
		);

	id_router_016 : component sopc_system_id_router_016
		port map (
			sink_ready         => sdram_0_avl_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sdram_0_avl_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sdram_0_avl_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sdram_0_avl_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sdram_0_avl_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => sdram_0_afi_clk_clk,                                                    --       clk.clk
			reset              => rst_controller_004_reset_out_reset,                                     -- clk_reset.reset
			src_ready          => id_router_016_src_ready,                                                --       src.ready
			src_valid          => id_router_016_src_valid,                                                --          .valid
			src_data           => id_router_016_src_data,                                                 --          .data
			src_channel        => id_router_016_src_channel,                                              --          .channel
			src_startofpacket  => id_router_016_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_016_src_endofpacket                                           --          .endofpacket
		);

	limiter : component sopc_system_limiter
		generic map (
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 88,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			MAX_OUTSTANDING_RESPONSES => 8,
			PIPELINED                 => 0,
			ST_DATA_W                 => 100,
			ST_CHANNEL_W              => 4,
			VALID_WIDTH               => 4,
			ENFORCE_ORDER             => 1,
			PREVENT_HAZARDS           => 0,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32
		)
		port map (
			clk                    => sdram_0_afi_clk_clk,                --       clk.clk
			reset                  => rst_controller_001_reset_out_reset, -- clk_reset.reset
			cmd_sink_ready         => addr_router_src_ready,              --  cmd_sink.ready
			cmd_sink_valid         => addr_router_src_valid,              --          .valid
			cmd_sink_data          => addr_router_src_data,               --          .data
			cmd_sink_channel       => addr_router_src_channel,            --          .channel
			cmd_sink_startofpacket => addr_router_src_startofpacket,      --          .startofpacket
			cmd_sink_endofpacket   => addr_router_src_endofpacket,        --          .endofpacket
			cmd_src_ready          => limiter_cmd_src_ready,              --   cmd_src.ready
			cmd_src_data           => limiter_cmd_src_data,               --          .data
			cmd_src_channel        => limiter_cmd_src_channel,            --          .channel
			cmd_src_startofpacket  => limiter_cmd_src_startofpacket,      --          .startofpacket
			cmd_src_endofpacket    => limiter_cmd_src_endofpacket,        --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_src_ready,             --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_src_valid,             --          .valid
			rsp_sink_channel       => rsp_xbar_mux_src_channel,           --          .channel
			rsp_sink_data          => rsp_xbar_mux_src_data,              --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_src_startofpacket,     --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_src_endofpacket,       --          .endofpacket
			rsp_src_ready          => limiter_rsp_src_ready,              --   rsp_src.ready
			rsp_src_valid          => limiter_rsp_src_valid,              --          .valid
			rsp_src_data           => limiter_rsp_src_data,               --          .data
			rsp_src_channel        => limiter_rsp_src_channel,            --          .channel
			rsp_src_startofpacket  => limiter_rsp_src_startofpacket,      --          .startofpacket
			rsp_src_endofpacket    => limiter_rsp_src_endofpacket,        --          .endofpacket
			cmd_src_valid          => limiter_cmd_valid_data              -- cmd_valid.data
		);

	limiter_001 : component sopc_system_limiter
		generic map (
			PKT_DEST_ID_H             => 89,
			PKT_DEST_ID_L             => 88,
			PKT_TRANS_POSTED          => 66,
			PKT_TRANS_WRITE           => 67,
			MAX_OUTSTANDING_RESPONSES => 8,
			PIPELINED                 => 0,
			ST_DATA_W                 => 100,
			ST_CHANNEL_W              => 4,
			VALID_WIDTH               => 4,
			ENFORCE_ORDER             => 1,
			PREVENT_HAZARDS           => 0,
			PKT_BYTE_CNT_H            => 73,
			PKT_BYTE_CNT_L            => 71,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32
		)
		port map (
			clk                    => sdram_0_afi_clk_clk,                --       clk.clk
			reset                  => rst_controller_001_reset_out_reset, -- clk_reset.reset
			cmd_sink_ready         => addr_router_001_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_001_src_valid,          --          .valid
			cmd_sink_data          => addr_router_001_src_data,           --          .data
			cmd_sink_channel       => addr_router_001_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_001_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_001_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_001_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_001_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_001_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_001_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_001_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_001_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_001_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_001_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_001_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_001_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_001_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_001_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_001_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_001_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_001_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_001_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_001_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_001_cmd_valid_data          -- cmd_valid.data
		);

	limiter_002 : component sopc_system_limiter_002
		generic map (
			PKT_DEST_ID_H             => 83,
			PKT_DEST_ID_L             => 81,
			PKT_TRANS_POSTED          => 60,
			PKT_TRANS_WRITE           => 61,
			MAX_OUTSTANDING_RESPONSES => 1,
			PIPELINED                 => 0,
			ST_DATA_W                 => 94,
			ST_CHANNEL_W              => 8,
			VALID_WIDTH               => 8,
			ENFORCE_ORDER             => 1,
			PREVENT_HAZARDS           => 0,
			PKT_BYTE_CNT_H            => 67,
			PKT_BYTE_CNT_L            => 65,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32
		)
		port map (
			clk                    => sdram_0_afi_half_clk_clk,           --       clk.clk
			reset                  => rst_controller_reset_out_reset,     -- clk_reset.reset
			cmd_sink_ready         => addr_router_007_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_007_src_valid,          --          .valid
			cmd_sink_data          => addr_router_007_src_data,           --          .data
			cmd_sink_channel       => addr_router_007_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_007_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_007_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_002_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_002_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_002_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_002_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_002_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_007_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_007_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_007_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_007_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_007_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_007_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_002_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_002_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_002_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_002_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_002_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_002_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_002_cmd_valid_data          -- cmd_valid.data
		);

	limiter_003 : component sopc_system_limiter_003
		generic map (
			PKT_DEST_ID_H             => 84,
			PKT_DEST_ID_L             => 84,
			PKT_TRANS_POSTED          => 65,
			PKT_TRANS_WRITE           => 66,
			MAX_OUTSTANDING_RESPONSES => 5,
			PIPELINED                 => 0,
			ST_DATA_W                 => 95,
			ST_CHANNEL_W              => 2,
			VALID_WIDTH               => 2,
			ENFORCE_ORDER             => 1,
			PREVENT_HAZARDS           => 0,
			PKT_BYTE_CNT_H            => 72,
			PKT_BYTE_CNT_L            => 70,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32
		)
		port map (
			clk                    => sdram_0_afi_half_clk_clk,           --       clk.clk
			reset                  => rst_controller_reset_out_reset,     -- clk_reset.reset
			cmd_sink_ready         => addr_router_008_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_008_src_valid,          --          .valid
			cmd_sink_data          => addr_router_008_src_data,           --          .data
			cmd_sink_channel       => addr_router_008_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_008_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_008_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_003_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_003_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_003_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_003_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_003_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_008_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_008_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_008_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_008_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_008_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_008_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_003_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_003_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_003_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_003_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_003_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_003_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_003_cmd_valid_data          -- cmd_valid.data
		);

	burst_adapter : component altera_merlin_burst_adapter
		generic map (
			PKT_ADDR_H                => 45,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 63,
			PKT_BYTE_CNT_H            => 54,
			PKT_BYTE_CNT_L            => 52,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 58,
			PKT_BURST_SIZE_L          => 56,
			PKT_BURST_TYPE_H          => 60,
			PKT_BURST_TYPE_L          => 59,
			PKT_BURSTWRAP_H           => 55,
			PKT_BURSTWRAP_L           => 55,
			PKT_TRANS_COMPRESSED_READ => 46,
			PKT_TRANS_WRITE           => 48,
			PKT_TRANS_READ            => 49,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 77,
			ST_CHANNEL_W              => 2,
			OUT_BYTE_CNT_H            => 53,
			OUT_BURSTWRAP_H           => 55,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 1,
			BURSTWRAP_CONST_VALUE     => 1
		)
		port map (
			clk                   => sdram_0_afi_half_clk_clk,            --       cr0.clk
			reset                 => rst_controller_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => width_adapter_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_src_data,              --          .data
			sink0_channel         => width_adapter_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_src_ready,             --          .ready
			source0_valid         => burst_adapter_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_source0_data,          --          .data
			source0_channel       => burst_adapter_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_source0_ready          --          .ready
		);

	burst_adapter_001 : component altera_merlin_burst_adapter
		generic map (
			PKT_ADDR_H                => 45,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 63,
			PKT_BYTE_CNT_H            => 54,
			PKT_BYTE_CNT_L            => 52,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 58,
			PKT_BURST_SIZE_L          => 56,
			PKT_BURST_TYPE_H          => 60,
			PKT_BURST_TYPE_L          => 59,
			PKT_BURSTWRAP_H           => 55,
			PKT_BURSTWRAP_L           => 55,
			PKT_TRANS_COMPRESSED_READ => 46,
			PKT_TRANS_WRITE           => 48,
			PKT_TRANS_READ            => 49,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 77,
			ST_CHANNEL_W              => 2,
			OUT_BYTE_CNT_H            => 53,
			OUT_BURSTWRAP_H           => 55,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 1,
			BURSTWRAP_CONST_VALUE     => 1
		)
		port map (
			clk                   => sdram_0_afi_half_clk_clk,                --       cr0.clk
			reset                 => rst_controller_reset_out_reset,          -- cr0_reset.reset
			sink0_valid           => width_adapter_002_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_002_src_data,              --          .data
			sink0_channel         => width_adapter_002_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_002_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_002_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_002_src_ready,             --          .ready
			source0_valid         => burst_adapter_001_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_001_source0_data,          --          .data
			source0_channel       => burst_adapter_001_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_001_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_001_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_001_source0_ready          --          .ready
		);

	rst_controller : component sopc_system_rst_controller
		generic map (
			NUM_RESET_INPUTS        => 3,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 1
		)
		port map (
			reset_in0  => linux_cpu_jtag_debug_module_reset_reset, -- reset_in0.reset
			reset_in1  => sdram_0_afi_reset_reset_ports_inv,       -- reset_in1.reset
			reset_in2  => clk_in_reset_reset_n_ports_inv,          -- reset_in2.reset
			clk        => sdram_0_afi_half_clk_clk,                --       clk.clk
			reset_out  => rst_controller_reset_out_reset,          -- reset_out.reset
			reset_req  => rst_controller_reset_out_reset_req,      --          .reset_req
			reset_in3  => '0',                                     -- (terminated)
			reset_in4  => '0',                                     -- (terminated)
			reset_in5  => '0',                                     -- (terminated)
			reset_in6  => '0',                                     -- (terminated)
			reset_in7  => '0',                                     -- (terminated)
			reset_in8  => '0',                                     -- (terminated)
			reset_in9  => '0',                                     -- (terminated)
			reset_in10 => '0',                                     -- (terminated)
			reset_in11 => '0',                                     -- (terminated)
			reset_in12 => '0',                                     -- (terminated)
			reset_in13 => '0',                                     -- (terminated)
			reset_in14 => '0',                                     -- (terminated)
			reset_in15 => '0'                                      -- (terminated)
		);

	rst_controller_001 : component sopc_system_rst_controller
		generic map (
			NUM_RESET_INPUTS        => 3,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 1
		)
		port map (
			reset_in0  => linux_cpu_jtag_debug_module_reset_reset, -- reset_in0.reset
			reset_in1  => sdram_0_afi_reset_reset_ports_inv,       -- reset_in1.reset
			reset_in2  => clk_in_reset_reset_n_ports_inv,          -- reset_in2.reset
			clk        => sdram_0_afi_clk_clk,                     --       clk.clk
			reset_out  => rst_controller_001_reset_out_reset,      -- reset_out.reset
			reset_req  => rst_controller_001_reset_out_reset_req,  --          .reset_req
			reset_in3  => '0',                                     -- (terminated)
			reset_in4  => '0',                                     -- (terminated)
			reset_in5  => '0',                                     -- (terminated)
			reset_in6  => '0',                                     -- (terminated)
			reset_in7  => '0',                                     -- (terminated)
			reset_in8  => '0',                                     -- (terminated)
			reset_in9  => '0',                                     -- (terminated)
			reset_in10 => '0',                                     -- (terminated)
			reset_in11 => '0',                                     -- (terminated)
			reset_in12 => '0',                                     -- (terminated)
			reset_in13 => '0',                                     -- (terminated)
			reset_in14 => '0',                                     -- (terminated)
			reset_in15 => '0'                                      -- (terminated)
		);

	rst_controller_002 : component sopc_system_rst_controller_002
		generic map (
			NUM_RESET_INPUTS        => 2,
			OUTPUT_RESET_SYNC_EDGES => "none",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => clk_in_reset_reset_n_ports_inv,          -- reset_in0.reset
			reset_in1  => linux_cpu_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk        => open,                                    --       clk.clk
			reset_out  => rst_controller_002_reset_out_reset,      -- reset_out.reset
			reset_req  => open,                                    -- (terminated)
			reset_in2  => '0',                                     -- (terminated)
			reset_in3  => '0',                                     -- (terminated)
			reset_in4  => '0',                                     -- (terminated)
			reset_in5  => '0',                                     -- (terminated)
			reset_in6  => '0',                                     -- (terminated)
			reset_in7  => '0',                                     -- (terminated)
			reset_in8  => '0',                                     -- (terminated)
			reset_in9  => '0',                                     -- (terminated)
			reset_in10 => '0',                                     -- (terminated)
			reset_in11 => '0',                                     -- (terminated)
			reset_in12 => '0',                                     -- (terminated)
			reset_in13 => '0',                                     -- (terminated)
			reset_in14 => '0',                                     -- (terminated)
			reset_in15 => '0'                                      -- (terminated)
		);

	rst_controller_003 : component sopc_system_rst_controller_003
		generic map (
			NUM_RESET_INPUTS        => 3,
			OUTPUT_RESET_SYNC_EDGES => "both",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => sdram_0_afi_reset_reset_ports_inv,       -- reset_in0.reset
			reset_in1  => clk_in_reset_reset_n_ports_inv,          -- reset_in1.reset
			reset_in2  => linux_cpu_jtag_debug_module_reset_reset, -- reset_in2.reset
			clk        => sdram_0_afi_half_clk_clk,                --       clk.clk
			reset_out  => rst_controller_003_reset_out_reset,      -- reset_out.reset
			reset_req  => open,                                    -- (terminated)
			reset_in3  => '0',                                     -- (terminated)
			reset_in4  => '0',                                     -- (terminated)
			reset_in5  => '0',                                     -- (terminated)
			reset_in6  => '0',                                     -- (terminated)
			reset_in7  => '0',                                     -- (terminated)
			reset_in8  => '0',                                     -- (terminated)
			reset_in9  => '0',                                     -- (terminated)
			reset_in10 => '0',                                     -- (terminated)
			reset_in11 => '0',                                     -- (terminated)
			reset_in12 => '0',                                     -- (terminated)
			reset_in13 => '0',                                     -- (terminated)
			reset_in14 => '0',                                     -- (terminated)
			reset_in15 => '0'                                      -- (terminated)
		);

	rst_controller_004 : component sopc_system_rst_controller_004
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => sdram_0_afi_reset_reset_ports_inv,  -- reset_in0.reset
			clk        => sdram_0_afi_clk_clk,                --       clk.clk
			reset_out  => rst_controller_004_reset_out_reset, -- reset_out.reset
			reset_req  => open,                               -- (terminated)
			reset_in1  => '0',                                -- (terminated)
			reset_in2  => '0',                                -- (terminated)
			reset_in3  => '0',                                -- (terminated)
			reset_in4  => '0',                                -- (terminated)
			reset_in5  => '0',                                -- (terminated)
			reset_in6  => '0',                                -- (terminated)
			reset_in7  => '0',                                -- (terminated)
			reset_in8  => '0',                                -- (terminated)
			reset_in9  => '0',                                -- (terminated)
			reset_in10 => '0',                                -- (terminated)
			reset_in11 => '0',                                -- (terminated)
			reset_in12 => '0',                                -- (terminated)
			reset_in13 => '0',                                -- (terminated)
			reset_in14 => '0',                                -- (terminated)
			reset_in15 => '0'                                 -- (terminated)
		);

	cmd_xbar_demux : component sopc_system_cmd_xbar_demux
		port map (
			clk                => sdram_0_afi_clk_clk,                --        clk.clk
			reset              => rst_controller_001_reset_out_reset, --  clk_reset.reset
			sink_ready         => limiter_cmd_src_ready,              --       sink.ready
			sink_channel       => limiter_cmd_src_channel,            --           .channel
			sink_data          => limiter_cmd_src_data,               --           .data
			sink_startofpacket => limiter_cmd_src_startofpacket,      --           .startofpacket
			sink_endofpacket   => limiter_cmd_src_endofpacket,        --           .endofpacket
			sink_valid         => limiter_cmd_valid_data,             -- sink_valid.data
			src0_ready         => cmd_xbar_demux_src0_ready,          --       src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,          --           .valid
			src0_data          => cmd_xbar_demux_src0_data,           --           .data
			src0_channel       => cmd_xbar_demux_src0_channel,        --           .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket,  --           .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,    --           .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,          --       src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,          --           .valid
			src1_data          => cmd_xbar_demux_src1_data,           --           .data
			src1_channel       => cmd_xbar_demux_src1_channel,        --           .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket,  --           .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket,    --           .endofpacket
			src2_ready         => cmd_xbar_demux_src2_ready,          --       src2.ready
			src2_valid         => cmd_xbar_demux_src2_valid,          --           .valid
			src2_data          => cmd_xbar_demux_src2_data,           --           .data
			src2_channel       => cmd_xbar_demux_src2_channel,        --           .channel
			src2_startofpacket => cmd_xbar_demux_src2_startofpacket,  --           .startofpacket
			src2_endofpacket   => cmd_xbar_demux_src2_endofpacket,    --           .endofpacket
			src3_ready         => cmd_xbar_demux_src3_ready,          --       src3.ready
			src3_valid         => cmd_xbar_demux_src3_valid,          --           .valid
			src3_data          => cmd_xbar_demux_src3_data,           --           .data
			src3_channel       => cmd_xbar_demux_src3_channel,        --           .channel
			src3_startofpacket => cmd_xbar_demux_src3_startofpacket,  --           .startofpacket
			src3_endofpacket   => cmd_xbar_demux_src3_endofpacket     --           .endofpacket
		);

	cmd_xbar_demux_001 : component sopc_system_cmd_xbar_demux_001
		port map (
			clk                => sdram_0_afi_clk_clk,                   --        clk.clk
			reset              => rst_controller_001_reset_out_reset,    --  clk_reset.reset
			sink_ready         => limiter_001_cmd_src_ready,             --       sink.ready
			sink_channel       => limiter_001_cmd_src_channel,           --           .channel
			sink_data          => limiter_001_cmd_src_data,              --           .data
			sink_startofpacket => limiter_001_cmd_src_startofpacket,     --           .startofpacket
			sink_endofpacket   => limiter_001_cmd_src_endofpacket,       --           .endofpacket
			sink_valid         => limiter_001_cmd_valid_data,            -- sink_valid.data
			src0_ready         => cmd_xbar_demux_001_src0_ready,         --       src0.ready
			src0_valid         => cmd_xbar_demux_001_src0_valid,         --           .valid
			src0_data          => cmd_xbar_demux_001_src0_data,          --           .data
			src0_channel       => cmd_xbar_demux_001_src0_channel,       --           .channel
			src0_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --           .startofpacket
			src0_endofpacket   => cmd_xbar_demux_001_src0_endofpacket,   --           .endofpacket
			src1_ready         => cmd_xbar_demux_001_src1_ready,         --       src1.ready
			src1_valid         => cmd_xbar_demux_001_src1_valid,         --           .valid
			src1_data          => cmd_xbar_demux_001_src1_data,          --           .data
			src1_channel       => cmd_xbar_demux_001_src1_channel,       --           .channel
			src1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --           .startofpacket
			src1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket,   --           .endofpacket
			src2_ready         => cmd_xbar_demux_001_src2_ready,         --       src2.ready
			src2_valid         => cmd_xbar_demux_001_src2_valid,         --           .valid
			src2_data          => cmd_xbar_demux_001_src2_data,          --           .data
			src2_channel       => cmd_xbar_demux_001_src2_channel,       --           .channel
			src2_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --           .startofpacket
			src2_endofpacket   => cmd_xbar_demux_001_src2_endofpacket    --           .endofpacket
		);

	cmd_xbar_mux : component sopc_system_cmd_xbar_mux
		port map (
			clk                 => sdram_0_afi_clk_clk,                   --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component sopc_system_cmd_xbar_mux
		port map (
			clk                 => sdram_0_afi_clk_clk,                   --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_003 : component sopc_system_cmd_xbar_mux
		port map (
			clk                 => sdram_0_afi_clk_clk,                   --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_003_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_003_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_003_src_data,             --          .data
			src_channel         => cmd_xbar_mux_003_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_003_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_003_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src3_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src3_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src3_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src3_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src3_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src3_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src2_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src2_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src2_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src2_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src2_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component sopc_system_rsp_xbar_demux
		port map (
			clk                => sdram_0_afi_clk_clk,                --       clk.clk
			reset              => rst_controller_001_reset_out_reset, -- clk_reset.reset
			sink_ready         => id_router_src_ready,                --      sink.ready
			sink_channel       => id_router_src_channel,              --          .channel
			sink_data          => id_router_src_data,                 --          .data
			sink_startofpacket => id_router_src_startofpacket,        --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,          --          .endofpacket
			sink_valid(0)      => id_router_src_valid,                --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,          --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,          --          .valid
			src0_data          => rsp_xbar_demux_src0_data,           --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,        --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket,  --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,    --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,          --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,          --          .valid
			src1_data          => rsp_xbar_demux_src1_data,           --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,        --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket,  --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket     --          .endofpacket
		);

	rsp_xbar_demux_001 : component sopc_system_rsp_xbar_demux
		port map (
			clk                => sdram_0_afi_clk_clk,                   --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_001_src_ready,               --      sink.ready
			sink_channel       => id_router_001_src_channel,             --          .channel
			sink_data          => id_router_001_src_data,                --          .data
			sink_startofpacket => id_router_001_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_001_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_001_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component sopc_system_rsp_xbar_demux_002
		port map (
			clk                => sdram_0_afi_clk_clk,                   --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component sopc_system_rsp_xbar_demux
		port map (
			clk                => sdram_0_afi_clk_clk,                   --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_003_src_ready,               --      sink.ready
			sink_channel       => id_router_003_src_channel,             --          .channel
			sink_data          => id_router_003_src_data,                --          .data
			sink_startofpacket => id_router_003_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_003_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_003_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_003_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_003_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_003_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_003_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_003_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component sopc_system_rsp_xbar_mux
		port map (
			clk                 => sdram_0_afi_clk_clk,                   --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready         => rsp_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			sink3_data          => rsp_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket   => rsp_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component sopc_system_rsp_xbar_mux_001
		port map (
			clk                 => sdram_0_afi_clk_clk,                   --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data            => rsp_xbar_mux_001_src_data,             --          .data
			src_channel         => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_003_src1_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_003_src1_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_003_src1_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_003_src1_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_003_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_002 : component sopc_system_cmd_xbar_demux_002
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_002_src_ready,             --      sink.ready
			sink_channel       => addr_router_002_src_channel,           --          .channel
			sink_data          => addr_router_002_src_data,              --          .data
			sink_startofpacket => addr_router_002_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_002_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_002_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_002_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_003 : component sopc_system_cmd_xbar_demux_002
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_003_src_ready,             --      sink.ready
			sink_channel       => addr_router_003_src_channel,           --          .channel
			sink_data          => addr_router_003_src_data,              --          .data
			sink_startofpacket => addr_router_003_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_003_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_003_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_003_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_004 : component sopc_system_cmd_xbar_demux_002
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_004_src_ready,             --      sink.ready
			sink_channel       => addr_router_004_src_channel,           --          .channel
			sink_data          => addr_router_004_src_data,              --          .data
			sink_startofpacket => addr_router_004_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_004_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_004_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_004_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_004_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_005 : component sopc_system_cmd_xbar_demux_002
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_005_src_ready,             --      sink.ready
			sink_channel       => addr_router_005_src_channel,           --          .channel
			sink_data          => addr_router_005_src_data,              --          .data
			sink_startofpacket => addr_router_005_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_005_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_005_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_005_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_005_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_004 : component sopc_system_cmd_xbar_mux_004
		port map (
			clk                 => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_004_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_004_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_004_src_data,             --          .data
			src_channel         => cmd_xbar_mux_004_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_004_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_004_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_002_src0_ready,         --     sink0.ready
			sink0_valid         => cmd_xbar_demux_002_src0_valid,         --          .valid
			sink0_channel       => cmd_xbar_demux_002_src0_channel,       --          .channel
			sink0_data          => cmd_xbar_demux_002_src0_data,          --          .data
			sink0_startofpacket => cmd_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink1_ready         => cmd_xbar_demux_003_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_003_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_003_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_003_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			sink2_ready         => cmd_xbar_demux_004_src0_ready,         --     sink2.ready
			sink2_valid         => cmd_xbar_demux_004_src0_valid,         --          .valid
			sink2_channel       => cmd_xbar_demux_004_src0_channel,       --          .channel
			sink2_data          => cmd_xbar_demux_004_src0_data,          --          .data
			sink2_startofpacket => cmd_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink2_endofpacket   => cmd_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			sink3_ready         => cmd_xbar_demux_005_src0_ready,         --     sink3.ready
			sink3_valid         => cmd_xbar_demux_005_src0_valid,         --          .valid
			sink3_channel       => cmd_xbar_demux_005_src0_channel,       --          .channel
			sink3_data          => cmd_xbar_demux_005_src0_data,          --          .data
			sink3_startofpacket => cmd_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink3_endofpacket   => cmd_xbar_demux_005_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component sopc_system_rsp_xbar_demux_004
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_004_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_004_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_004_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_004_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_004_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_004_src1_endofpacket,   --          .endofpacket
			src2_ready         => rsp_xbar_demux_004_src2_ready,         --      src2.ready
			src2_valid         => rsp_xbar_demux_004_src2_valid,         --          .valid
			src2_data          => rsp_xbar_demux_004_src2_data,          --          .data
			src2_channel       => rsp_xbar_demux_004_src2_channel,       --          .channel
			src2_startofpacket => rsp_xbar_demux_004_src2_startofpacket, --          .startofpacket
			src2_endofpacket   => rsp_xbar_demux_004_src2_endofpacket,   --          .endofpacket
			src3_ready         => rsp_xbar_demux_004_src3_ready,         --      src3.ready
			src3_valid         => rsp_xbar_demux_004_src3_valid,         --          .valid
			src3_data          => rsp_xbar_demux_004_src3_data,          --          .data
			src3_channel       => rsp_xbar_demux_004_src3_channel,       --          .channel
			src3_startofpacket => rsp_xbar_demux_004_src3_startofpacket, --          .startofpacket
			src3_endofpacket   => rsp_xbar_demux_004_src3_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_006 : component sopc_system_cmd_xbar_demux_006
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_006_src_ready,             --      sink.ready
			sink_channel       => addr_router_006_src_channel,           --          .channel
			sink_data          => addr_router_006_src_data,              --          .data
			sink_startofpacket => addr_router_006_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_006_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_006_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_006_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_007 : component sopc_system_cmd_xbar_demux_007
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --        clk.clk
			reset              => rst_controller_reset_out_reset,        --  clk_reset.reset
			sink_ready         => limiter_002_cmd_src_ready,             --       sink.ready
			sink_channel       => limiter_002_cmd_src_channel,           --           .channel
			sink_data          => limiter_002_cmd_src_data,              --           .data
			sink_startofpacket => limiter_002_cmd_src_startofpacket,     --           .startofpacket
			sink_endofpacket   => limiter_002_cmd_src_endofpacket,       --           .endofpacket
			sink_valid         => limiter_002_cmd_valid_data,            -- sink_valid.data
			src0_ready         => cmd_xbar_demux_007_src0_ready,         --       src0.ready
			src0_valid         => cmd_xbar_demux_007_src0_valid,         --           .valid
			src0_data          => cmd_xbar_demux_007_src0_data,          --           .data
			src0_channel       => cmd_xbar_demux_007_src0_channel,       --           .channel
			src0_startofpacket => cmd_xbar_demux_007_src0_startofpacket, --           .startofpacket
			src0_endofpacket   => cmd_xbar_demux_007_src0_endofpacket,   --           .endofpacket
			src1_ready         => cmd_xbar_demux_007_src1_ready,         --       src1.ready
			src1_valid         => cmd_xbar_demux_007_src1_valid,         --           .valid
			src1_data          => cmd_xbar_demux_007_src1_data,          --           .data
			src1_channel       => cmd_xbar_demux_007_src1_channel,       --           .channel
			src1_startofpacket => cmd_xbar_demux_007_src1_startofpacket, --           .startofpacket
			src1_endofpacket   => cmd_xbar_demux_007_src1_endofpacket,   --           .endofpacket
			src2_ready         => cmd_xbar_demux_007_src2_ready,         --       src2.ready
			src2_valid         => cmd_xbar_demux_007_src2_valid,         --           .valid
			src2_data          => cmd_xbar_demux_007_src2_data,          --           .data
			src2_channel       => cmd_xbar_demux_007_src2_channel,       --           .channel
			src2_startofpacket => cmd_xbar_demux_007_src2_startofpacket, --           .startofpacket
			src2_endofpacket   => cmd_xbar_demux_007_src2_endofpacket,   --           .endofpacket
			src3_ready         => cmd_xbar_demux_007_src3_ready,         --       src3.ready
			src3_valid         => cmd_xbar_demux_007_src3_valid,         --           .valid
			src3_data          => cmd_xbar_demux_007_src3_data,          --           .data
			src3_channel       => cmd_xbar_demux_007_src3_channel,       --           .channel
			src3_startofpacket => cmd_xbar_demux_007_src3_startofpacket, --           .startofpacket
			src3_endofpacket   => cmd_xbar_demux_007_src3_endofpacket,   --           .endofpacket
			src4_ready         => cmd_xbar_demux_007_src4_ready,         --       src4.ready
			src4_valid         => cmd_xbar_demux_007_src4_valid,         --           .valid
			src4_data          => cmd_xbar_demux_007_src4_data,          --           .data
			src4_channel       => cmd_xbar_demux_007_src4_channel,       --           .channel
			src4_startofpacket => cmd_xbar_demux_007_src4_startofpacket, --           .startofpacket
			src4_endofpacket   => cmd_xbar_demux_007_src4_endofpacket,   --           .endofpacket
			src5_ready         => cmd_xbar_demux_007_src5_ready,         --       src5.ready
			src5_valid         => cmd_xbar_demux_007_src5_valid,         --           .valid
			src5_data          => cmd_xbar_demux_007_src5_data,          --           .data
			src5_channel       => cmd_xbar_demux_007_src5_channel,       --           .channel
			src5_startofpacket => cmd_xbar_demux_007_src5_startofpacket, --           .startofpacket
			src5_endofpacket   => cmd_xbar_demux_007_src5_endofpacket,   --           .endofpacket
			src6_ready         => cmd_xbar_demux_007_src6_ready,         --       src6.ready
			src6_valid         => cmd_xbar_demux_007_src6_valid,         --           .valid
			src6_data          => cmd_xbar_demux_007_src6_data,          --           .data
			src6_channel       => cmd_xbar_demux_007_src6_channel,       --           .channel
			src6_startofpacket => cmd_xbar_demux_007_src6_startofpacket, --           .startofpacket
			src6_endofpacket   => cmd_xbar_demux_007_src6_endofpacket,   --           .endofpacket
			src7_ready         => cmd_xbar_demux_007_src7_ready,         --       src7.ready
			src7_valid         => cmd_xbar_demux_007_src7_valid,         --           .valid
			src7_data          => cmd_xbar_demux_007_src7_data,          --           .data
			src7_channel       => cmd_xbar_demux_007_src7_channel,       --           .channel
			src7_startofpacket => cmd_xbar_demux_007_src7_startofpacket, --           .startofpacket
			src7_endofpacket   => cmd_xbar_demux_007_src7_endofpacket    --           .endofpacket
		);

	cmd_xbar_mux_005 : component sopc_system_cmd_xbar_mux_005
		port map (
			clk                 => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_005_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_005_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_005_src_data,             --          .data
			src_channel         => cmd_xbar_mux_005_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_005_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_005_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_006_src0_ready,         --     sink0.ready
			sink0_valid         => cmd_xbar_demux_006_src0_valid,         --          .valid
			sink0_channel       => cmd_xbar_demux_006_src0_channel,       --          .channel
			sink0_data          => cmd_xbar_demux_006_src0_data,          --          .data
			sink0_startofpacket => cmd_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			sink1_ready         => cmd_xbar_demux_007_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_007_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_007_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_007_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component sopc_system_rsp_xbar_demux_005
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_005_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_005_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_005_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_005_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_005_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_005_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component sopc_system_cmd_xbar_demux_006
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component sopc_system_cmd_xbar_demux_006
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_008 : component sopc_system_cmd_xbar_demux_006
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_008_src_ready,               --      sink.ready
			sink_channel       => id_router_008_src_channel,             --          .channel
			sink_data          => id_router_008_src_data,                --          .data
			sink_startofpacket => id_router_008_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_008_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_008_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_008_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_008_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_008_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_009 : component sopc_system_cmd_xbar_demux_006
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_009_src_ready,               --      sink.ready
			sink_channel       => id_router_009_src_channel,             --          .channel
			sink_data          => id_router_009_src_data,                --          .data
			sink_startofpacket => id_router_009_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_009_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_009_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_009_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_010 : component sopc_system_cmd_xbar_demux_006
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_010_src_ready,               --      sink.ready
			sink_channel       => id_router_010_src_channel,             --          .channel
			sink_data          => id_router_010_src_data,                --          .data
			sink_startofpacket => id_router_010_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_010_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_010_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_010_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_010_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_010_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_011 : component sopc_system_cmd_xbar_demux_006
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_011_src_ready,               --      sink.ready
			sink_channel       => id_router_011_src_channel,             --          .channel
			sink_data          => id_router_011_src_data,                --          .data
			sink_startofpacket => id_router_011_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_011_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_011_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_011_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_011_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_011_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_012 : component sopc_system_cmd_xbar_demux_006
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_012_src_ready,               --      sink.ready
			sink_channel       => id_router_012_src_channel,             --          .channel
			sink_data          => id_router_012_src_data,                --          .data
			sink_startofpacket => id_router_012_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_012_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_012_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_012_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_012_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_012_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_007 : component sopc_system_rsp_xbar_mux_007
		port map (
			clk                 => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_007_src_ready,            --       src.ready
			src_valid           => rsp_xbar_mux_007_src_valid,            --          .valid
			src_data            => rsp_xbar_mux_007_src_data,             --          .data
			src_channel         => rsp_xbar_mux_007_src_channel,          --          .channel
			src_startofpacket   => rsp_xbar_mux_007_src_startofpacket,    --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_007_src_endofpacket,      --          .endofpacket
			sink0_ready         => rsp_xbar_demux_005_src1_ready,         --     sink0.ready
			sink0_valid         => rsp_xbar_demux_005_src1_valid,         --          .valid
			sink0_channel       => rsp_xbar_demux_005_src1_channel,       --          .channel
			sink0_data          => rsp_xbar_demux_005_src1_data,          --          .data
			sink0_startofpacket => rsp_xbar_demux_005_src1_startofpacket, --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_005_src1_endofpacket,   --          .endofpacket
			sink1_ready         => rsp_xbar_demux_006_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_006_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_007_src0_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_007_src0_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			sink3_ready         => rsp_xbar_demux_008_src0_ready,         --     sink3.ready
			sink3_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			sink3_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			sink3_data          => rsp_xbar_demux_008_src0_data,          --          .data
			sink3_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			sink3_endofpacket   => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			sink4_ready         => rsp_xbar_demux_009_src0_ready,         --     sink4.ready
			sink4_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			sink4_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			sink4_data          => rsp_xbar_demux_009_src0_data,          --          .data
			sink4_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			sink4_endofpacket   => rsp_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			sink5_ready         => rsp_xbar_demux_010_src0_ready,         --     sink5.ready
			sink5_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			sink5_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			sink5_data          => rsp_xbar_demux_010_src0_data,          --          .data
			sink5_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			sink5_endofpacket   => rsp_xbar_demux_010_src0_endofpacket,   --          .endofpacket
			sink6_ready         => rsp_xbar_demux_011_src0_ready,         --     sink6.ready
			sink6_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			sink6_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			sink6_data          => rsp_xbar_demux_011_src0_data,          --          .data
			sink6_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			sink6_endofpacket   => rsp_xbar_demux_011_src0_endofpacket,   --          .endofpacket
			sink7_ready         => rsp_xbar_demux_012_src0_ready,         --     sink7.ready
			sink7_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			sink7_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			sink7_data          => rsp_xbar_demux_012_src0_data,          --          .data
			sink7_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			sink7_endofpacket   => rsp_xbar_demux_012_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_008 : component sopc_system_cmd_xbar_demux_008
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --        clk.clk
			reset              => rst_controller_reset_out_reset,        --  clk_reset.reset
			sink_ready         => limiter_003_cmd_src_ready,             --       sink.ready
			sink_channel       => limiter_003_cmd_src_channel,           --           .channel
			sink_data          => limiter_003_cmd_src_data,              --           .data
			sink_startofpacket => limiter_003_cmd_src_startofpacket,     --           .startofpacket
			sink_endofpacket   => limiter_003_cmd_src_endofpacket,       --           .endofpacket
			sink_valid         => limiter_003_cmd_valid_data,            -- sink_valid.data
			src0_ready         => cmd_xbar_demux_008_src0_ready,         --       src0.ready
			src0_valid         => cmd_xbar_demux_008_src0_valid,         --           .valid
			src0_data          => cmd_xbar_demux_008_src0_data,          --           .data
			src0_channel       => cmd_xbar_demux_008_src0_channel,       --           .channel
			src0_startofpacket => cmd_xbar_demux_008_src0_startofpacket, --           .startofpacket
			src0_endofpacket   => cmd_xbar_demux_008_src0_endofpacket,   --           .endofpacket
			src1_ready         => cmd_xbar_demux_008_src1_ready,         --       src1.ready
			src1_valid         => cmd_xbar_demux_008_src1_valid,         --           .valid
			src1_data          => cmd_xbar_demux_008_src1_data,          --           .data
			src1_channel       => cmd_xbar_demux_008_src1_channel,       --           .channel
			src1_startofpacket => cmd_xbar_demux_008_src1_startofpacket, --           .startofpacket
			src1_endofpacket   => cmd_xbar_demux_008_src1_endofpacket    --           .endofpacket
		);

	rsp_xbar_demux_013 : component sopc_system_rsp_xbar_demux_013
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => width_adapter_001_src_ready,           --      sink.ready
			sink_channel       => width_adapter_001_src_channel,         --          .channel
			sink_data          => width_adapter_001_src_data,            --          .data
			sink_startofpacket => width_adapter_001_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_001_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_001_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_013_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_013_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_013_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_014 : component sopc_system_rsp_xbar_demux_013
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => width_adapter_003_src_ready,           --      sink.ready
			sink_channel       => width_adapter_003_src_channel,         --          .channel
			sink_data          => width_adapter_003_src_data,            --          .data
			sink_startofpacket => width_adapter_003_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_003_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_003_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_014_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_014_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_014_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_008 : component sopc_system_rsp_xbar_mux_008
		port map (
			clk                 => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_008_src_ready,            --       src.ready
			src_valid           => rsp_xbar_mux_008_src_valid,            --          .valid
			src_data            => rsp_xbar_mux_008_src_data,             --          .data
			src_channel         => rsp_xbar_mux_008_src_channel,          --          .channel
			src_startofpacket   => rsp_xbar_mux_008_src_startofpacket,    --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_008_src_endofpacket,      --          .endofpacket
			sink0_ready         => rsp_xbar_demux_013_src0_ready,         --     sink0.ready
			sink0_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			sink0_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			sink0_data          => rsp_xbar_demux_013_src0_data,          --          .data
			sink0_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_013_src0_endofpacket,   --          .endofpacket
			sink1_ready         => rsp_xbar_demux_014_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_014_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_014_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_009 : component sopc_system_cmd_xbar_demux_009
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_009_src_ready,             --      sink.ready
			sink_channel       => addr_router_009_src_channel,           --          .channel
			sink_data          => addr_router_009_src_data,              --          .data
			sink_startofpacket => addr_router_009_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_009_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_009_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_009_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_010 : component sopc_system_cmd_xbar_demux_009
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_010_src_ready,             --      sink.ready
			sink_channel       => addr_router_010_src_channel,           --          .channel
			sink_data          => addr_router_010_src_data,              --          .data
			sink_startofpacket => addr_router_010_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_010_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_010_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_010_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_010_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_010_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_010_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_010_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_010_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_015 : component sopc_system_cmd_xbar_mux_015
		port map (
			clk                 => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_015_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_015_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_015_src_data,             --          .data
			src_channel         => cmd_xbar_mux_015_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_015_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_015_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_009_src0_ready,         --     sink0.ready
			sink0_valid         => cmd_xbar_demux_009_src0_valid,         --          .valid
			sink0_channel       => cmd_xbar_demux_009_src0_channel,       --          .channel
			sink0_data          => cmd_xbar_demux_009_src0_data,          --          .data
			sink0_startofpacket => cmd_xbar_demux_009_src0_startofpacket, --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			sink1_ready         => cmd_xbar_demux_010_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_010_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_010_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_010_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_010_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_010_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_015 : component sopc_system_rsp_xbar_demux_015
		port map (
			clk                => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_015_src_ready,               --      sink.ready
			sink_channel       => id_router_015_src_channel,             --          .channel
			sink_data          => id_router_015_src_data,                --          .data
			sink_startofpacket => id_router_015_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_015_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_015_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_015_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_015_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_015_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_015_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_015_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_015_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_015_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_015_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_015_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_015_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_015_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_015_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_011 : component sopc_system_cmd_xbar_demux_011
		port map (
			clk                => sdram_0_afi_clk_clk,                   --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => addr_router_011_src_ready,             --      sink.ready
			sink_channel       => addr_router_011_src_channel,           --          .channel
			sink_data          => addr_router_011_src_data,              --          .data
			sink_startofpacket => addr_router_011_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_011_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_011_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_011_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_011_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_011_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_011_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_011_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_011_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_012 : component sopc_system_cmd_xbar_demux_011
		port map (
			clk                => sdram_0_afi_clk_clk,                   --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => addr_router_012_src_ready,             --      sink.ready
			sink_channel       => addr_router_012_src_channel,           --          .channel
			sink_data          => addr_router_012_src_data,              --          .data
			sink_startofpacket => addr_router_012_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_012_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_012_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_012_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_012_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_012_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_012_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_012_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_012_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_016 : component sopc_system_cmd_xbar_mux_016
		port map (
			clk                 => sdram_0_afi_clk_clk,                   --       clk.clk
			reset               => rst_controller_004_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_016_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_016_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_016_src_data,             --          .data
			src_channel         => cmd_xbar_mux_016_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_016_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_016_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_011_src0_ready,         --     sink0.ready
			sink0_valid         => cmd_xbar_demux_011_src0_valid,         --          .valid
			sink0_channel       => cmd_xbar_demux_011_src0_channel,       --          .channel
			sink0_data          => cmd_xbar_demux_011_src0_data,          --          .data
			sink0_startofpacket => cmd_xbar_demux_011_src0_startofpacket, --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_011_src0_endofpacket,   --          .endofpacket
			sink1_ready         => cmd_xbar_demux_012_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_012_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_012_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_012_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_012_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_012_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_016 : component sopc_system_rsp_xbar_demux_016
		port map (
			clk                => sdram_0_afi_clk_clk,                   --       clk.clk
			reset              => rst_controller_004_reset_out_reset,    -- clk_reset.reset
			sink_ready         => width_adapter_005_src_ready,           --      sink.ready
			sink_channel       => width_adapter_005_src_channel,         --          .channel
			sink_data          => width_adapter_005_src_data,            --          .data
			sink_startofpacket => width_adapter_005_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_005_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_005_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_016_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_016_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_016_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_016_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_016_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_016_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_016_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_016_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_016_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_016_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_016_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_016_src1_endofpacket    --          .endofpacket
		);

	width_adapter : component sopc_system_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 63,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 72,
			IN_PKT_BYTE_CNT_L             => 70,
			IN_PKT_TRANS_COMPRESSED_READ  => 64,
			IN_PKT_BURSTWRAP_H            => 73,
			IN_PKT_BURSTWRAP_L            => 73,
			IN_PKT_BURST_SIZE_H           => 76,
			IN_PKT_BURST_SIZE_L           => 74,
			IN_PKT_RESPONSE_STATUS_H      => 94,
			IN_PKT_RESPONSE_STATUS_L      => 93,
			IN_PKT_TRANS_EXCLUSIVE        => 69,
			IN_PKT_BURST_TYPE_H           => 78,
			IN_PKT_BURST_TYPE_L           => 77,
			IN_ST_DATA_W                  => 95,
			OUT_PKT_ADDR_H                => 45,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 54,
			OUT_PKT_BYTE_CNT_L            => 52,
			OUT_PKT_TRANS_COMPRESSED_READ => 46,
			OUT_PKT_BURST_SIZE_H          => 58,
			OUT_PKT_BURST_SIZE_L          => 56,
			OUT_PKT_RESPONSE_STATUS_H     => 76,
			OUT_PKT_RESPONSE_STATUS_L     => 75,
			OUT_PKT_TRANS_EXCLUSIVE       => 51,
			OUT_PKT_BURST_TYPE_H          => 60,
			OUT_PKT_BURST_TYPE_L          => 59,
			OUT_ST_DATA_W                 => 77,
			ST_CHANNEL_W                  => 2,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => cmd_xbar_demux_008_src0_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_008_src0_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_008_src0_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_008_src0_ready,         --          .ready
			in_data              => cmd_xbar_demux_008_src0_data,          --          .data
			out_endofpacket      => width_adapter_src_endofpacket,         --       src.endofpacket
			out_data             => width_adapter_src_data,                --          .data
			out_channel          => width_adapter_src_channel,             --          .channel
			out_valid            => width_adapter_src_valid,               --          .valid
			out_ready            => width_adapter_src_ready,               --          .ready
			out_startofpacket    => width_adapter_src_startofpacket,       --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_001 : component sopc_system_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 45,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 54,
			IN_PKT_BYTE_CNT_L             => 52,
			IN_PKT_TRANS_COMPRESSED_READ  => 46,
			IN_PKT_BURSTWRAP_H            => 55,
			IN_PKT_BURSTWRAP_L            => 55,
			IN_PKT_BURST_SIZE_H           => 58,
			IN_PKT_BURST_SIZE_L           => 56,
			IN_PKT_RESPONSE_STATUS_H      => 76,
			IN_PKT_RESPONSE_STATUS_L      => 75,
			IN_PKT_TRANS_EXCLUSIVE        => 51,
			IN_PKT_BURST_TYPE_H           => 60,
			IN_PKT_BURST_TYPE_L           => 59,
			IN_ST_DATA_W                  => 77,
			OUT_PKT_ADDR_H                => 63,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 72,
			OUT_PKT_BYTE_CNT_L            => 70,
			OUT_PKT_TRANS_COMPRESSED_READ => 64,
			OUT_PKT_BURST_SIZE_H          => 76,
			OUT_PKT_BURST_SIZE_L          => 74,
			OUT_PKT_RESPONSE_STATUS_H     => 94,
			OUT_PKT_RESPONSE_STATUS_L     => 93,
			OUT_PKT_TRANS_EXCLUSIVE       => 69,
			OUT_PKT_BURST_TYPE_H          => 78,
			OUT_PKT_BURST_TYPE_L          => 77,
			OUT_ST_DATA_W                 => 95,
			ST_CHANNEL_W                  => 2,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => sdram_0_afi_half_clk_clk,            --       clk.clk
			reset                => rst_controller_reset_out_reset,      -- clk_reset.reset
			in_valid             => id_router_013_src_valid,             --      sink.valid
			in_channel           => id_router_013_src_channel,           --          .channel
			in_startofpacket     => id_router_013_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_013_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_013_src_ready,             --          .ready
			in_data              => id_router_013_src_data,              --          .data
			out_endofpacket      => width_adapter_001_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_001_src_data,          --          .data
			out_channel          => width_adapter_001_src_channel,       --          .channel
			out_valid            => width_adapter_001_src_valid,         --          .valid
			out_ready            => width_adapter_001_src_ready,         --          .ready
			out_startofpacket    => width_adapter_001_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_002 : component sopc_system_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 63,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 72,
			IN_PKT_BYTE_CNT_L             => 70,
			IN_PKT_TRANS_COMPRESSED_READ  => 64,
			IN_PKT_BURSTWRAP_H            => 73,
			IN_PKT_BURSTWRAP_L            => 73,
			IN_PKT_BURST_SIZE_H           => 76,
			IN_PKT_BURST_SIZE_L           => 74,
			IN_PKT_RESPONSE_STATUS_H      => 94,
			IN_PKT_RESPONSE_STATUS_L      => 93,
			IN_PKT_TRANS_EXCLUSIVE        => 69,
			IN_PKT_BURST_TYPE_H           => 78,
			IN_PKT_BURST_TYPE_L           => 77,
			IN_ST_DATA_W                  => 95,
			OUT_PKT_ADDR_H                => 45,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 54,
			OUT_PKT_BYTE_CNT_L            => 52,
			OUT_PKT_TRANS_COMPRESSED_READ => 46,
			OUT_PKT_BURST_SIZE_H          => 58,
			OUT_PKT_BURST_SIZE_L          => 56,
			OUT_PKT_RESPONSE_STATUS_H     => 76,
			OUT_PKT_RESPONSE_STATUS_L     => 75,
			OUT_PKT_TRANS_EXCLUSIVE       => 51,
			OUT_PKT_BURST_TYPE_H          => 60,
			OUT_PKT_BURST_TYPE_L          => 59,
			OUT_ST_DATA_W                 => 77,
			ST_CHANNEL_W                  => 2,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => sdram_0_afi_half_clk_clk,              --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			in_valid             => cmd_xbar_demux_008_src1_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_008_src1_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_008_src1_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_008_src1_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_008_src1_ready,         --          .ready
			in_data              => cmd_xbar_demux_008_src1_data,          --          .data
			out_endofpacket      => width_adapter_002_src_endofpacket,     --       src.endofpacket
			out_data             => width_adapter_002_src_data,            --          .data
			out_channel          => width_adapter_002_src_channel,         --          .channel
			out_valid            => width_adapter_002_src_valid,           --          .valid
			out_ready            => width_adapter_002_src_ready,           --          .ready
			out_startofpacket    => width_adapter_002_src_startofpacket,   --          .startofpacket
			in_command_size_data => "000"                                  -- (terminated)
		);

	width_adapter_003 : component sopc_system_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 45,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 54,
			IN_PKT_BYTE_CNT_L             => 52,
			IN_PKT_TRANS_COMPRESSED_READ  => 46,
			IN_PKT_BURSTWRAP_H            => 55,
			IN_PKT_BURSTWRAP_L            => 55,
			IN_PKT_BURST_SIZE_H           => 58,
			IN_PKT_BURST_SIZE_L           => 56,
			IN_PKT_RESPONSE_STATUS_H      => 76,
			IN_PKT_RESPONSE_STATUS_L      => 75,
			IN_PKT_TRANS_EXCLUSIVE        => 51,
			IN_PKT_BURST_TYPE_H           => 60,
			IN_PKT_BURST_TYPE_L           => 59,
			IN_ST_DATA_W                  => 77,
			OUT_PKT_ADDR_H                => 63,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 72,
			OUT_PKT_BYTE_CNT_L            => 70,
			OUT_PKT_TRANS_COMPRESSED_READ => 64,
			OUT_PKT_BURST_SIZE_H          => 76,
			OUT_PKT_BURST_SIZE_L          => 74,
			OUT_PKT_RESPONSE_STATUS_H     => 94,
			OUT_PKT_RESPONSE_STATUS_L     => 93,
			OUT_PKT_TRANS_EXCLUSIVE       => 69,
			OUT_PKT_BURST_TYPE_H          => 78,
			OUT_PKT_BURST_TYPE_L          => 77,
			OUT_ST_DATA_W                 => 95,
			ST_CHANNEL_W                  => 2,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => sdram_0_afi_half_clk_clk,            --       clk.clk
			reset                => rst_controller_reset_out_reset,      -- clk_reset.reset
			in_valid             => id_router_014_src_valid,             --      sink.valid
			in_channel           => id_router_014_src_channel,           --          .channel
			in_startofpacket     => id_router_014_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_014_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_014_src_ready,             --          .ready
			in_data              => id_router_014_src_data,              --          .data
			out_endofpacket      => width_adapter_003_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_003_src_data,          --          .data
			out_channel          => width_adapter_003_src_channel,       --          .channel
			out_valid            => width_adapter_003_src_valid,         --          .valid
			out_ready            => width_adapter_003_src_ready,         --          .ready
			out_startofpacket    => width_adapter_003_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_004 : component sopc_system_width_adapter_004
		generic map (
			IN_PKT_ADDR_H                 => 62,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 74,
			IN_PKT_BYTE_CNT_L             => 69,
			IN_PKT_TRANS_COMPRESSED_READ  => 63,
			IN_PKT_BURSTWRAP_H            => 75,
			IN_PKT_BURSTWRAP_L            => 75,
			IN_PKT_BURST_SIZE_H           => 78,
			IN_PKT_BURST_SIZE_L           => 76,
			IN_PKT_RESPONSE_STATUS_H      => 96,
			IN_PKT_RESPONSE_STATUS_L      => 95,
			IN_PKT_TRANS_EXCLUSIVE        => 68,
			IN_PKT_BURST_TYPE_H           => 80,
			IN_PKT_BURST_TYPE_L           => 79,
			IN_ST_DATA_W                  => 97,
			OUT_PKT_ADDR_H                => 98,
			OUT_PKT_ADDR_L                => 72,
			OUT_PKT_DATA_H                => 63,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 71,
			OUT_PKT_BYTEEN_L              => 64,
			OUT_PKT_BYTE_CNT_H            => 110,
			OUT_PKT_BYTE_CNT_L            => 105,
			OUT_PKT_TRANS_COMPRESSED_READ => 99,
			OUT_PKT_BURST_SIZE_H          => 114,
			OUT_PKT_BURST_SIZE_L          => 112,
			OUT_PKT_RESPONSE_STATUS_H     => 132,
			OUT_PKT_RESPONSE_STATUS_L     => 131,
			OUT_PKT_TRANS_EXCLUSIVE       => 104,
			OUT_PKT_BURST_TYPE_H          => 116,
			OUT_PKT_BURST_TYPE_L          => 115,
			OUT_ST_DATA_W                 => 133,
			ST_CHANNEL_W                  => 2,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => sdram_0_afi_clk_clk,                 --       clk.clk
			reset                => rst_controller_004_reset_out_reset,  -- clk_reset.reset
			in_valid             => cmd_xbar_mux_016_src_valid,          --      sink.valid
			in_channel           => cmd_xbar_mux_016_src_channel,        --          .channel
			in_startofpacket     => cmd_xbar_mux_016_src_startofpacket,  --          .startofpacket
			in_endofpacket       => cmd_xbar_mux_016_src_endofpacket,    --          .endofpacket
			in_ready             => cmd_xbar_mux_016_src_ready,          --          .ready
			in_data              => cmd_xbar_mux_016_src_data,           --          .data
			out_endofpacket      => width_adapter_004_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_004_src_data,          --          .data
			out_channel          => width_adapter_004_src_channel,       --          .channel
			out_valid            => width_adapter_004_src_valid,         --          .valid
			out_ready            => width_adapter_004_src_ready,         --          .ready
			out_startofpacket    => width_adapter_004_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_005 : component sopc_system_width_adapter_005
		generic map (
			IN_PKT_ADDR_H                 => 98,
			IN_PKT_ADDR_L                 => 72,
			IN_PKT_DATA_H                 => 63,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 71,
			IN_PKT_BYTEEN_L               => 64,
			IN_PKT_BYTE_CNT_H             => 110,
			IN_PKT_BYTE_CNT_L             => 105,
			IN_PKT_TRANS_COMPRESSED_READ  => 99,
			IN_PKT_BURSTWRAP_H            => 111,
			IN_PKT_BURSTWRAP_L            => 111,
			IN_PKT_BURST_SIZE_H           => 114,
			IN_PKT_BURST_SIZE_L           => 112,
			IN_PKT_RESPONSE_STATUS_H      => 132,
			IN_PKT_RESPONSE_STATUS_L      => 131,
			IN_PKT_TRANS_EXCLUSIVE        => 104,
			IN_PKT_BURST_TYPE_H           => 116,
			IN_PKT_BURST_TYPE_L           => 115,
			IN_ST_DATA_W                  => 133,
			OUT_PKT_ADDR_H                => 62,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 74,
			OUT_PKT_BYTE_CNT_L            => 69,
			OUT_PKT_TRANS_COMPRESSED_READ => 63,
			OUT_PKT_BURST_SIZE_H          => 78,
			OUT_PKT_BURST_SIZE_L          => 76,
			OUT_PKT_RESPONSE_STATUS_H     => 96,
			OUT_PKT_RESPONSE_STATUS_L     => 95,
			OUT_PKT_TRANS_EXCLUSIVE       => 68,
			OUT_PKT_BURST_TYPE_H          => 80,
			OUT_PKT_BURST_TYPE_L          => 79,
			OUT_ST_DATA_W                 => 97,
			ST_CHANNEL_W                  => 2,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => sdram_0_afi_clk_clk,                 --       clk.clk
			reset                => rst_controller_004_reset_out_reset,  -- clk_reset.reset
			in_valid             => id_router_016_src_valid,             --      sink.valid
			in_channel           => id_router_016_src_channel,           --          .channel
			in_startofpacket     => id_router_016_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_016_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_016_src_ready,             --          .ready
			in_data              => id_router_016_src_data,              --          .data
			out_endofpacket      => width_adapter_005_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_005_src_data,          --          .data
			out_channel          => width_adapter_005_src_channel,       --          .channel
			out_valid            => width_adapter_005_src_valid,         --          .valid
			out_ready            => width_adapter_005_src_ready,         --          .ready
			out_startofpacket    => width_adapter_005_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	irq_mapper : component sopc_system_irq_mapper
		port map (
			clk           => sdram_0_afi_clk_clk,                --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			sender_irq    => linux_cpu_d_irq_irq                 --    sender.irq
		);

	irq_synchronizer : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => sdram_0_afi_half_clk_clk,           --       receiver_clk.clk
			sender_clk     => sdram_0_afi_clk_clk,                --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_receiver_irq,      --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver0_irq            --             sender.irq
		);

	irq_synchronizer_001 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => sdram_0_afi_half_clk_clk,           --       receiver_clk.clk
			sender_clk     => sdram_0_afi_clk_clk,                --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_001_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver1_irq            --             sender.irq
		);

	irq_synchronizer_002 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => sdram_0_afi_half_clk_clk,           --       receiver_clk.clk
			sender_clk     => sdram_0_afi_clk_clk,                --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_002_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver2_irq            --             sender.irq
		);

	irq_synchronizer_003 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => sdram_0_afi_half_clk_clk,           --       receiver_clk.clk
			sender_clk     => sdram_0_afi_clk_clk,                --         sender_clk.clk
			receiver_reset => rst_controller_reset_out_reset,     -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_003_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver3_irq            --             sender.irq
		);

	irq_synchronizer_004 : component altera_irq_clock_crosser
		generic map (
			IRQ_WIDTH => 1
		)
		port map (
			receiver_clk   => sdram_0_afi_half_clk_clk,           --       receiver_clk.clk
			sender_clk     => sdram_0_afi_clk_clk,                --         sender_clk.clk
			receiver_reset => rst_controller_003_reset_out_reset, -- receiver_clk_reset.reset
			sender_reset   => rst_controller_001_reset_out_reset, --   sender_clk_reset.reset
			receiver_irq   => irq_synchronizer_004_receiver_irq,  --           receiver.irq
			sender_irq(0)  => irq_mapper_receiver4_irq            --             sender.irq
		);

	avalon_st_adapter : component sopc_system_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 6,
			inUseEmptyPort  => 1,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 2,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 6,
			outUseEmptyPort => 1,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => sdram_0_afi_half_clk_clk,              -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,        -- in_rst_0.reset
			in_0_ready          => tse_mac_receive_ready,                 --     in_0.ready
			in_0_valid          => tse_mac_receive_valid,                 --         .valid
			in_0_data           => tse_mac_receive_data,                  --         .data
			in_0_startofpacket  => tse_mac_receive_startofpacket,         --         .startofpacket
			in_0_endofpacket    => tse_mac_receive_endofpacket,           --         .endofpacket
			in_0_empty          => tse_mac_receive_empty,                 --         .empty
			in_0_error          => tse_mac_receive_error,                 --         .error
			out_0_ready         => avalon_st_adapter_out_0_ready,         --    out_0.ready
			out_0_valid         => avalon_st_adapter_out_0_valid,         --         .valid
			out_0_data          => avalon_st_adapter_out_0_data,          --         .data
			out_0_startofpacket => avalon_st_adapter_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_out_0_endofpacket,   --         .endofpacket
			out_0_empty         => avalon_st_adapter_out_0_empty,         --         .empty
			out_0_error         => avalon_st_adapter_out_0_error          --         .error
		);

	clk_in_reset_reset_n_ports_inv <= not clk_in_reset_reset_n;

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	linux_timer_1ms_s1_translator_avalon_anti_slave_0_write_ports_inv <= not linux_timer_1ms_s1_translator_avalon_anti_slave_0_write;

	sdram_0_avl_translator_avalon_anti_slave_0_inv <= not sdram_0_avl_waitrequest;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	sdram_0_afi_reset_reset_ports_inv <= not sdram_0_afi_reset_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

end architecture rtl; -- of sopc_system
